******************************************************************
** Silicon Creations Confidential
** LVS Netlist for PLLTS40GFRAC - Version v3d53
** This netlist is intended to be used for layout comparison (LVS)
** Not intended for SPICE simulation
**
**
**

.subckt nmoscap_18 PLUS MINUS lr=1u wr=1u m=1
.ends

.subckt PLLTS40GFRAC BYPASS CLKSSCG DACPD DSMPD FBDIV[0] FBDIV[10] FBDIV[11]
+ FBDIV[1] FBDIV[2] FBDIV[3] FBDIV[4] FBDIV[5] FBDIV[6] FBDIV[7] FBDIV[8]
+ FBDIV[9] FOUT1PH0 FOUT1PH180 FOUT1PH270 FOUT1PH90 FOUT2 FOUT3 FOUT4
+ FOUT4PHASEPD FOUTPOSTDIV FOUTPOSTDIVPD FOUTVCO FOUTVCOPD FRAC[0] FRAC[10]
+ FRAC[11] FRAC[12] FRAC[13] FRAC[14] FRAC[15] FRAC[16] FRAC[17] FRAC[18]
+ FRAC[19] FRAC[1] FRAC[20] FRAC[21] FRAC[22] FRAC[23] FRAC[2] FRAC[3] FRAC[4]
+ FRAC[5] FRAC[6] FRAC[7] FRAC[8] FRAC[9] FREF LOCK PD POSTDIV1[0] POSTDIV1[1]
+ POSTDIV1[2] POSTDIV2[0] POSTDIV2[1] POSTDIV2[2] REFDIV[0] REFDIV[1] REFDIV[2]
+ REFDIV[3] REFDIV[4] REFDIV[5] VDDHV VDDPOST VDDREF VSS
m0 5490 5313 2 VSS nch_18 l=0.28u w=0.44u
m1 5067 5316 5490 VSS nch_18 l=0.28u w=0.44u
m2 5725 5313 5067 VSS nch_18 l=0.28u w=0.44u
m3 5786 5316 5725 VSS nch_18 l=0.28u w=0.44u
m4 VSS 4948 4795 VSS nch_18 l=0.55u w=0.44u
m5 4796 4795 VSS VSS nch_18 l=0.55u w=0.44u
m6 VSS 4869 4864 VSS nch_18 l=0.55u w=0.44u
m7 4865 4859 VSS VSS nch_18 l=0.55u w=0.44u
m8 VSS 4949 4869 VSS nch_18 l=0.55u w=0.44u
m9 4869 4795 VSS VSS nch_18 l=0.55u w=0.44u
m10 4861 4795 2 VSS nch_18 l=0.55u w=2.08u
m11 VSS 4869 4861 VSS nch_18 l=0.55u w=2.08u
m12 4862 4795 VSS VSS nch_18 l=0.55u w=2.08u
m13 2 4869 4862 VSS nch_18 l=0.55u w=2.08u
m14 VSS 4940 4859 VSS nch_18 l=0.55u w=5.44u
m15 4946 4943 VSS VSS nch_18 l=0.55u w=5.44u
m16 VSS 4961 4954 VSS nch_18 l=0.55u w=5.44u
m17 4948 4964 VSS VSS nch_18 l=0.55u w=5.44u
m18 VSS 4979 4971 VSS nch_18 l=0.55u w=5.44u
m19 4949 4983 VSS VSS nch_18 l=0.55u w=5.44u
m20 72213 4994 VSS VSS nch_18 l=0.65u w=1.3u
m21 72214 4994 VSS VSS nch_18 l=0.65u w=1.3u
m22 72215 4994 VSS VSS nch_18 l=0.65u w=1.3u
m23 72216 4994 VSS VSS nch_18 l=0.65u w=1.3u
m24 5000 5858 4994 VSS nch_18 l=0.55u w=0.65u
m25 VSS 4992 4996 VSS nch_18 l=0.55u w=0.44u
m26 5016 5040 4992 VSS nch_18 l=0.55u w=2u
m27 4994 5858 5000 VSS nch_18 l=0.55u w=0.65u
m28 72223 4994 72213 VSS nch_18 l=0.65u w=1.3u
m29 72224 4994 72214 VSS nch_18 l=0.65u w=1.3u
m30 72225 4994 72215 VSS nch_18 l=0.65u w=1.3u
m31 72226 4994 72216 VSS nch_18 l=0.65u w=1.3u
m32 5020 4996 VSS VSS nch_18 l=0.55u w=0.44u
m33 5020 4996 VSS VSS nch_18 l=0.55u w=0.44u
m34 5000 5858 4994 VSS nch_18 l=0.55u w=0.65u
m35 72230 4994 72223 VSS nch_18 l=0.65u w=1.3u
m36 72231 4994 72224 VSS nch_18 l=0.65u w=1.3u
m37 72232 4994 72225 VSS nch_18 l=0.65u w=1.3u
m38 72233 4994 72226 VSS nch_18 l=0.65u w=1.3u
m39 5040 5040 VDDREF VSS nch_18 l=0.55u w=2u
m40 VSS 4996 5020 VSS nch_18 l=0.55u w=0.44u
m41 VSS 4996 5020 VSS nch_18 l=0.55u w=0.44u
m42 4994 5858 5000 VSS nch_18 l=0.55u w=0.65u
m43 5000 4994 72230 VSS nch_18 l=0.65u w=1.3u
m44 5000 4994 72231 VSS nch_18 l=0.65u w=1.3u
m45 5000 4994 72232 VSS nch_18 l=0.65u w=1.3u
m46 5000 4994 72233 VSS nch_18 l=0.65u w=1.3u
m47 5048 5072 VSS VSS nch_18 l=0.55u w=0.44u
m48 5048 5072 VSS VSS nch_18 l=0.55u w=0.44u
m49 VDDREF 5040 5040 VSS nch_18 l=0.55u w=2u
m50 VSS 5072 5048 VSS nch_18 l=0.55u w=0.44u
m51 VSS 5072 5048 VSS nch_18 l=0.55u w=0.44u
m52 5068 5040 5050 VSS nch_18 l=0.55u w=2u
m53 72254 4994 VSS VSS nch_18 l=0.65u w=1.3u
m54 72255 4994 VSS VSS nch_18 l=0.65u w=1.3u
m55 72256 4994 VSS VSS nch_18 l=0.65u w=1.3u
m56 72257 4994 VSS VSS nch_18 l=0.65u w=1.3u
m57 5072 5068 VSS VSS nch_18 l=0.55u w=0.44u
m58 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m59 5091 VDDHV VSS VSS nch_18 l=5u w=0.44u
m60 5091 VDDHV 4992 VSS nch_18 l=5u w=0.44u
m61 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m62 72266 4994 72254 VSS nch_18 l=0.65u w=1.3u
m63 72267 4994 72255 VSS nch_18 l=0.65u w=1.3u
m64 72268 4994 72256 VSS nch_18 l=0.65u w=1.3u
m65 72269 4994 72257 VSS nch_18 l=0.65u w=1.3u
m66 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m67 VSS 5093 5097 VSS nch_18 l=0.55u w=0.44u
m68 72274 4994 72266 VSS nch_18 l=0.65u w=1.3u
m69 72275 4994 72267 VSS nch_18 l=0.65u w=1.3u
m70 72276 4994 72268 VSS nch_18 l=0.65u w=1.3u
m71 72277 4994 72269 VSS nch_18 l=0.65u w=1.3u
m72 5116 5139 5093 VSS nch_18 l=0.55u w=2u
m73 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m74 5131 5097 VSS VSS nch_18 l=0.55u w=0.44u
m75 5131 5097 VSS VSS nch_18 l=0.55u w=0.44u
m76 5086 4994 72274 VSS nch_18 l=0.65u w=1.3u
m77 5086 4994 72275 VSS nch_18 l=0.65u w=1.3u
m78 5086 4994 72276 VSS nch_18 l=0.65u w=1.3u
m79 5086 4994 72277 VSS nch_18 l=0.65u w=1.3u
m80 5139 5139 VDDREF VSS nch_18 l=0.55u w=2u
m81 VSS 5097 5131 VSS nch_18 l=0.55u w=0.44u
m82 VSS 5097 5131 VSS nch_18 l=0.55u w=0.44u
m83 5158 5183 VSS VSS nch_18 l=0.55u w=0.44u
m84 5158 5183 VSS VSS nch_18 l=0.55u w=0.44u
m85 VDDREF 5139 5139 VSS nch_18 l=0.55u w=2u
m86 72292 4994 VSS VSS nch_18 l=0.65u w=1.3u
m87 72293 4994 VSS VSS nch_18 l=0.65u w=1.3u
m88 72294 4994 VSS VSS nch_18 l=0.65u w=1.3u
m89 72295 4994 VSS VSS nch_18 l=0.65u w=1.3u
m90 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m91 VSS 5183 5158 VSS nch_18 l=0.55u w=0.44u
m92 VSS 5183 5158 VSS nch_18 l=0.55u w=0.44u
m93 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m94 72299 4994 72292 VSS nch_18 l=0.65u w=1.3u
m95 72300 4994 72293 VSS nch_18 l=0.65u w=1.3u
m96 72301 4994 72294 VSS nch_18 l=0.65u w=1.3u
m97 72302 4994 72295 VSS nch_18 l=0.65u w=1.3u
m98 5178 5139 5159 VSS nch_18 l=0.55u w=2u
m99 5183 5178 VSS VSS nch_18 l=0.55u w=0.44u
m100 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m101 5190 VDDHV VSS VSS nch_18 l=5u w=0.44u
m102 5190 VDDHV 5093 VSS nch_18 l=5u w=0.44u
m103 72308 4994 72299 VSS nch_18 l=0.65u w=1.3u
m104 72309 4994 72300 VSS nch_18 l=0.65u w=1.3u
m105 72310 4994 72301 VSS nch_18 l=0.65u w=1.3u
m106 72311 4994 72302 VSS nch_18 l=0.65u w=1.3u
m107 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m108 5086 4994 72308 VSS nch_18 l=0.65u w=1.3u
m109 5086 4994 72309 VSS nch_18 l=0.65u w=1.3u
m110 5086 4994 72310 VSS nch_18 l=0.65u w=1.3u
m111 5086 4994 72311 VSS nch_18 l=0.65u w=1.3u
m112 VSS 5048 5205 VSS nch_18 l=0.55u w=0.44u
m113 VSS 5205 5206 VSS nch_18 l=0.55u w=2u
m114 5231 5020 VSS VSS nch_18 l=0.55u w=0.44u
m115 5230 5234 VSS VSS nch_18 l=0.55u w=2u
m116 5234 5205 VSS VSS nch_18 l=0.55u w=0.44u
m117 72341 4994 VSS VSS nch_18 l=0.65u w=1.3u
m118 72342 4994 VSS VSS nch_18 l=0.65u w=1.3u
m119 72343 4994 VSS VSS nch_18 l=0.65u w=1.3u
m120 72344 4994 VSS VSS nch_18 l=0.65u w=1.3u
m121 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m122 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m123 72355 4994 72341 VSS nch_18 l=0.65u w=1.3u
m124 72356 4994 72342 VSS nch_18 l=0.65u w=1.3u
m125 72357 4994 72343 VSS nch_18 l=0.65u w=1.3u
m126 72358 4994 72344 VSS nch_18 l=0.65u w=1.3u
m127 VSS 5273 5249 VSS nch_18 l=0.55u w=0.44u
m128 VSS 5131 5250 VSS nch_18 l=0.55u w=0.44u
m129 VSS 5249 5251 VSS nch_18 l=0.55u w=2u
m130 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m131 72367 4994 72355 VSS nch_18 l=0.65u w=1.3u
m132 72368 4994 72356 VSS nch_18 l=0.65u w=1.3u
m133 72369 4994 72357 VSS nch_18 l=0.65u w=1.3u
m134 72370 4994 72358 VSS nch_18 l=0.65u w=1.3u
m135 5273 5158 VSS VSS nch_18 l=0.55u w=0.44u
m136 5274 5273 VSS VSS nch_18 l=0.55u w=2u
m137 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m138 5086 4994 72367 VSS nch_18 l=0.65u w=1.3u
m139 5086 4994 72368 VSS nch_18 l=0.65u w=1.3u
m140 5086 4994 72369 VSS nch_18 l=0.65u w=1.3u
m141 5086 4994 72370 VSS nch_18 l=0.65u w=1.3u
m142 72404 4994 VSS VSS nch_18 l=0.65u w=1.3u
m143 72405 4994 VSS VSS nch_18 l=0.65u w=1.3u
m144 72406 4994 VSS VSS nch_18 l=0.65u w=1.3u
m145 72407 4994 VSS VSS nch_18 l=0.65u w=1.3u
m146 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m147 5312 5131 VSS VSS nch_18 l=0.55u w=0.44u
m148 5313 5312 VSS VSS nch_18 l=0.55u w=0.44u
m149 5314 5357 VSS VSS nch_18 l=0.55u w=0.44u
m150 5315 5158 VSS VSS nch_18 l=0.55u w=0.44u
m151 5316 5315 VSS VSS nch_18 l=0.55u w=0.44u
m152 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m153 72410 4994 72404 VSS nch_18 l=0.65u w=1.3u
m154 72411 4994 72405 VSS nch_18 l=0.65u w=1.3u
m155 72412 4994 72406 VSS nch_18 l=0.65u w=1.3u
m156 72413 4994 72407 VSS nch_18 l=0.65u w=1.3u
m157 VSS 5131 5312 VSS nch_18 l=0.55u w=0.44u
m158 VSS 5312 5313 VSS nch_18 l=0.55u w=0.44u
m159 VSS 5357 5314 VSS nch_18 l=0.55u w=0.44u
m160 VSS 5158 5315 VSS nch_18 l=0.55u w=0.44u
m161 VSS 5315 5316 VSS nch_18 l=0.55u w=0.44u
m162 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m163 5359 5020 VSS VSS nch_18 l=0.55u w=0.44u
m164 5357 5359 VSS VSS nch_18 l=0.55u w=0.44u
m165 5360 5356 VSS VSS nch_18 l=0.55u w=0.44u
m166 5358 5048 VSS VSS nch_18 l=0.55u w=0.44u
m167 5356 5358 VSS VSS nch_18 l=0.55u w=0.44u
m168 72416 4994 72410 VSS nch_18 l=0.65u w=1.3u
m169 72417 4994 72411 VSS nch_18 l=0.65u w=1.3u
m170 72418 4994 72412 VSS nch_18 l=0.65u w=1.3u
m171 72419 4994 72413 VSS nch_18 l=0.65u w=1.3u
m172 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m173 VSS 5020 5359 VSS nch_18 l=0.55u w=0.44u
m174 VSS 5359 5357 VSS nch_18 l=0.55u w=0.44u
m175 VSS 5356 5360 VSS nch_18 l=0.55u w=0.44u
m176 VSS 5048 5358 VSS nch_18 l=0.55u w=0.44u
m177 VSS 5358 5356 VSS nch_18 l=0.55u w=0.44u
m178 5086 4994 72416 VSS nch_18 l=0.65u w=1.3u
m179 5086 4994 72417 VSS nch_18 l=0.65u w=1.3u
m180 5086 4994 72418 VSS nch_18 l=0.65u w=1.3u
m181 5086 4994 72419 VSS nch_18 l=0.65u w=1.3u
m182 72447 4994 VSS VSS nch_18 l=0.65u w=1.3u
m183 72448 4994 VSS VSS nch_18 l=0.65u w=1.3u
m184 72449 4994 VSS VSS nch_18 l=0.65u w=1.3u
m185 72450 4994 VSS VSS nch_18 l=0.65u w=1.3u
m186 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m187 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m188 72504 4994 72447 VSS nch_18 l=0.65u w=1.3u
m189 72505 4994 72448 VSS nch_18 l=0.65u w=1.3u
m190 72506 4994 72449 VSS nch_18 l=0.65u w=1.3u
m191 72507 4994 72450 VSS nch_18 l=0.65u w=1.3u
m192 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m193 72508 4994 72504 VSS nch_18 l=0.65u w=1.3u
m194 72509 4994 72505 VSS nch_18 l=0.65u w=1.3u
m195 72510 4994 72506 VSS nch_18 l=0.65u w=1.3u
m196 72511 4994 72507 VSS nch_18 l=0.65u w=1.3u
m197 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m198 5086 4994 72508 VSS nch_18 l=0.65u w=1.3u
m199 5086 4994 72509 VSS nch_18 l=0.65u w=1.3u
m200 5086 4994 72510 VSS nch_18 l=0.65u w=1.3u
m201 5086 4994 72511 VSS nch_18 l=0.65u w=1.3u
m202 72561 5809 5489 VSS nch_18 l=0.65u w=1.3u
m203 72562 5809 5489 VSS nch_18 l=0.65u w=1.3u
m204 72563 5809 5489 VSS nch_18 l=0.65u w=1.3u
m205 72564 5809 5489 VSS nch_18 l=0.65u w=1.3u
m206 5489 5823 5490 VSS nch_18 l=0.55u w=0.65u
m207 72570 4994 VSS VSS nch_18 l=0.65u w=1.3u
m208 72571 4994 VSS VSS nch_18 l=0.65u w=1.3u
m209 72572 4994 VSS VSS nch_18 l=0.65u w=1.3u
m210 72573 4994 VSS VSS nch_18 l=0.65u w=1.3u
m211 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m212 5490 5823 5489 VSS nch_18 l=0.55u w=0.65u
m213 72576 5809 72561 VSS nch_18 l=0.65u w=1.3u
m214 72577 5809 72562 VSS nch_18 l=0.65u w=1.3u
m215 72578 5809 72563 VSS nch_18 l=0.65u w=1.3u
m216 72579 5809 72564 VSS nch_18 l=0.65u w=1.3u
m217 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m218 72589 4994 72570 VSS nch_18 l=0.65u w=1.3u
m219 72590 4994 72571 VSS nch_18 l=0.65u w=1.3u
m220 72591 4994 72572 VSS nch_18 l=0.65u w=1.3u
m221 72592 4994 72573 VSS nch_18 l=0.65u w=1.3u
m222 5489 5823 5490 VSS nch_18 l=0.55u w=0.65u
m223 72596 5809 72576 VSS nch_18 l=0.65u w=1.3u
m224 72597 5809 72577 VSS nch_18 l=0.65u w=1.3u
m225 72598 5809 72578 VSS nch_18 l=0.65u w=1.3u
m226 72599 5809 72579 VSS nch_18 l=0.65u w=1.3u
m227 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m228 72608 4994 72589 VSS nch_18 l=0.65u w=1.3u
m229 72609 4994 72590 VSS nch_18 l=0.65u w=1.3u
m230 72610 4994 72591 VSS nch_18 l=0.65u w=1.3u
m231 72611 4994 72592 VSS nch_18 l=0.65u w=1.3u
m232 5595 5595 VSS VSS nch_18 l=0.78u w=0.975u
m233 5490 5823 5489 VSS nch_18 l=0.55u w=0.65u
m234 VSS 5809 72596 VSS nch_18 l=0.65u w=1.3u
m235 VSS 5809 72597 VSS nch_18 l=0.65u w=1.3u
m236 VSS 5809 72598 VSS nch_18 l=0.65u w=1.3u
m237 VSS 5809 72599 VSS nch_18 l=0.65u w=1.3u
m238 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m239 5086 4994 72608 VSS nch_18 l=0.65u w=1.3u
m240 5086 4994 72609 VSS nch_18 l=0.65u w=1.3u
m241 5086 4994 72610 VSS nch_18 l=0.65u w=1.3u
m242 5086 4994 72611 VSS nch_18 l=0.65u w=1.3u
m243 VSS 5595 5595 VSS nch_18 l=0.78u w=0.975u
m244 72648 5809 5610 VSS nch_18 l=0.65u w=1.3u
m245 72649 5809 5610 VSS nch_18 l=0.65u w=1.3u
m246 72650 5809 5610 VSS nch_18 l=0.65u w=1.3u
m247 72651 5809 5610 VSS nch_18 l=0.65u w=1.3u
m248 5643 5595 VSS VSS nch_18 l=0.78u w=0.975u
m249 72662 4994 VSS VSS nch_18 l=0.65u w=1.3u
m250 72663 4994 VSS VSS nch_18 l=0.65u w=1.3u
m251 72664 4994 VSS VSS nch_18 l=0.65u w=1.3u
m252 72665 4994 VSS VSS nch_18 l=0.65u w=1.3u
m253 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m254 72675 5809 72648 VSS nch_18 l=0.65u w=1.3u
m255 72676 5809 72649 VSS nch_18 l=0.65u w=1.3u
m256 72677 5809 72650 VSS nch_18 l=0.65u w=1.3u
m257 72678 5809 72651 VSS nch_18 l=0.65u w=1.3u
m258 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m259 72691 4994 72662 VSS nch_18 l=0.65u w=1.3u
m260 72692 4994 72663 VSS nch_18 l=0.65u w=1.3u
m261 72693 4994 72664 VSS nch_18 l=0.65u w=1.3u
m262 72694 4994 72665 VSS nch_18 l=0.65u w=1.3u
m263 VSS 5595 5643 VSS nch_18 l=0.78u w=0.975u
m264 72700 5809 72675 VSS nch_18 l=0.65u w=1.3u
m265 72701 5809 72676 VSS nch_18 l=0.65u w=1.3u
m266 72702 5809 72677 VSS nch_18 l=0.65u w=1.3u
m267 72703 5809 72678 VSS nch_18 l=0.65u w=1.3u
m268 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m269 72715 4994 72691 VSS nch_18 l=0.65u w=1.3u
m270 72716 4994 72692 VSS nch_18 l=0.65u w=1.3u
m271 72717 4994 72693 VSS nch_18 l=0.65u w=1.3u
m272 72718 4994 72694 VSS nch_18 l=0.65u w=1.3u
m273 VSS 5809 72700 VSS nch_18 l=0.65u w=1.3u
m274 VSS 5809 72701 VSS nch_18 l=0.65u w=1.3u
m275 VSS 5809 72702 VSS nch_18 l=0.65u w=1.3u
m276 VSS 5809 72703 VSS nch_18 l=0.65u w=1.3u
m277 5595 5595 VSS VSS nch_18 l=0.78u w=0.975u
m278 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m279 5086 4994 72715 VSS nch_18 l=0.65u w=1.3u
m280 5086 4994 72716 VSS nch_18 l=0.65u w=1.3u
m281 5086 4994 72717 VSS nch_18 l=0.65u w=1.3u
m282 5086 4994 72718 VSS nch_18 l=0.65u w=1.3u
m283 VSS 5595 5595 VSS nch_18 l=0.78u w=0.975u
m284 72754 5809 5723 VSS nch_18 l=0.65u w=1.3u
m285 72755 5809 5723 VSS nch_18 l=0.65u w=1.3u
m286 72756 5809 5723 VSS nch_18 l=0.65u w=1.3u
m287 72757 5809 5723 VSS nch_18 l=0.65u w=1.3u
m288 5723 5823 5725 VSS nch_18 l=0.55u w=0.65u
m289 72769 4994 VSS VSS nch_18 l=0.65u w=1.3u
m290 72770 4994 VSS VSS nch_18 l=0.65u w=1.3u
m291 72771 4994 VSS VSS nch_18 l=0.65u w=1.3u
m292 72772 4994 VSS VSS nch_18 l=0.65u w=1.3u
m293 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m294 5643 5595 VSS VSS nch_18 l=0.78u w=0.975u
m295 5725 5823 5723 VSS nch_18 l=0.55u w=0.65u
m296 72776 5809 72754 VSS nch_18 l=0.65u w=1.3u
m297 72777 5809 72755 VSS nch_18 l=0.65u w=1.3u
m298 72778 5809 72756 VSS nch_18 l=0.65u w=1.3u
m299 72779 5809 72757 VSS nch_18 l=0.65u w=1.3u
m300 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m301 72793 4994 72769 VSS nch_18 l=0.65u w=1.3u
m302 72794 4994 72770 VSS nch_18 l=0.65u w=1.3u
m303 72795 4994 72771 VSS nch_18 l=0.65u w=1.3u
m304 72796 4994 72772 VSS nch_18 l=0.65u w=1.3u
m305 5723 5823 5725 VSS nch_18 l=0.55u w=0.65u
m306 72804 5809 72776 VSS nch_18 l=0.65u w=1.3u
m307 72805 5809 72777 VSS nch_18 l=0.65u w=1.3u
m308 72806 5809 72778 VSS nch_18 l=0.65u w=1.3u
m309 72807 5809 72779 VSS nch_18 l=0.65u w=1.3u
m310 VSS 5595 5643 VSS nch_18 l=0.78u w=0.975u
m311 5086 5858 5067 VSS nch_18 l=0.55u w=0.65u
m312 72817 4994 72793 VSS nch_18 l=0.65u w=1.3u
m313 72818 4994 72794 VSS nch_18 l=0.65u w=1.3u
m314 72819 4994 72795 VSS nch_18 l=0.65u w=1.3u
m315 72820 4994 72796 VSS nch_18 l=0.65u w=1.3u
m316 5725 5823 5723 VSS nch_18 l=0.55u w=0.65u
m317 VSS 5809 72804 VSS nch_18 l=0.65u w=1.3u
m318 VSS 5809 72805 VSS nch_18 l=0.65u w=1.3u
m319 VSS 5809 72806 VSS nch_18 l=0.65u w=1.3u
m320 VSS 5809 72807 VSS nch_18 l=0.65u w=1.3u
m321 5067 5858 5086 VSS nch_18 l=0.55u w=0.65u
m322 5086 4994 72817 VSS nch_18 l=0.65u w=1.3u
m323 5086 4994 72818 VSS nch_18 l=0.65u w=1.3u
m324 5086 4994 72819 VSS nch_18 l=0.65u w=1.3u
m325 5086 4994 72820 VSS nch_18 l=0.65u w=1.3u
m326 72869 5823 5791 VSS nch_18 l=0.65u w=1.3u
m327 72870 5823 5791 VSS nch_18 l=0.65u w=1.3u
m328 72871 5823 5791 VSS nch_18 l=0.65u w=1.3u
m329 72872 5823 5791 VSS nch_18 l=0.65u w=1.3u
m330 72891 4994 VSS VSS nch_18 l=0.65u w=1.3u
m331 72892 4994 VSS VSS nch_18 l=0.65u w=1.3u
m332 72893 4994 VSS VSS nch_18 l=0.65u w=1.3u
m333 72894 4994 VSS VSS nch_18 l=0.65u w=1.3u
m334 5800 5858 5786 VSS nch_18 l=0.55u w=0.65u
m335 72900 5823 72869 VSS nch_18 l=0.65u w=1.3u
m336 72901 5823 72870 VSS nch_18 l=0.65u w=1.3u
m337 72902 5823 72871 VSS nch_18 l=0.65u w=1.3u
m338 72903 5823 72872 VSS nch_18 l=0.65u w=1.3u
m339 5786 5858 5800 VSS nch_18 l=0.55u w=0.65u
m340 72922 4994 72891 VSS nch_18 l=0.65u w=1.3u
m341 72923 4994 72892 VSS nch_18 l=0.65u w=1.3u
m342 72924 4994 72893 VSS nch_18 l=0.65u w=1.3u
m343 72925 4994 72894 VSS nch_18 l=0.65u w=1.3u
m344 72930 5823 72900 VSS nch_18 l=0.65u w=1.3u
m345 72931 5823 72901 VSS nch_18 l=0.65u w=1.3u
m346 72932 5823 72902 VSS nch_18 l=0.65u w=1.3u
m347 72933 5823 72903 VSS nch_18 l=0.65u w=1.3u
m348 5800 5858 5786 VSS nch_18 l=0.55u w=0.65u
m349 72949 4994 72922 VSS nch_18 l=0.65u w=1.3u
m350 72950 4994 72923 VSS nch_18 l=0.65u w=1.3u
m351 72951 4994 72924 VSS nch_18 l=0.65u w=1.3u
m352 72952 4994 72925 VSS nch_18 l=0.65u w=1.3u
m353 5823 5823 72930 VSS nch_18 l=0.65u w=1.3u
m354 5823 5823 72931 VSS nch_18 l=0.65u w=1.3u
m355 VSS 5823 72932 VSS nch_18 l=0.65u w=1.3u
m356 VSS 5823 72933 VSS nch_18 l=0.65u w=1.3u
m357 5786 5858 5800 VSS nch_18 l=0.55u w=0.65u
m358 5800 4994 72949 VSS nch_18 l=0.65u w=1.3u
m359 5800 4994 72950 VSS nch_18 l=0.65u w=1.3u
m360 5800 4994 72951 VSS nch_18 l=0.65u w=1.3u
m361 5800 4994 72952 VSS nch_18 l=0.65u w=1.3u
m362 72994 5809 5828 VSS nch_18 l=0.65u w=1.3u
m363 72995 5809 5828 VSS nch_18 l=0.65u w=1.3u
m364 72996 5809 5828 VSS nch_18 l=0.65u w=1.3u
m365 72997 5809 5828 VSS nch_18 l=0.65u w=1.3u
m366 5828 5823 5809 VSS nch_18 l=0.55u w=0.65u
m367 73006 4994 VSS VSS nch_18 l=0.65u w=1.3u
m368 73007 4994 VSS VSS nch_18 l=0.65u w=1.3u
m369 73008 4994 VSS VSS nch_18 l=0.65u w=1.3u
m370 73009 4994 VSS VSS nch_18 l=0.65u w=1.3u
m371 5800 5858 5786 VSS nch_18 l=0.55u w=0.65u
m372 5809 5823 5828 VSS nch_18 l=0.55u w=0.65u
m373 73013 5809 72994 VSS nch_18 l=0.65u w=1.3u
m374 73014 5809 72995 VSS nch_18 l=0.65u w=1.3u
m375 73015 5809 72996 VSS nch_18 l=0.65u w=1.3u
m376 73016 5809 72997 VSS nch_18 l=0.65u w=1.3u
m377 5786 5858 5800 VSS nch_18 l=0.55u w=0.65u
m378 73028 4994 73006 VSS nch_18 l=0.65u w=1.3u
m379 73029 4994 73007 VSS nch_18 l=0.65u w=1.3u
m380 73030 4994 73008 VSS nch_18 l=0.65u w=1.3u
m381 73031 4994 73009 VSS nch_18 l=0.65u w=1.3u
m382 5828 5823 5809 VSS nch_18 l=0.55u w=0.65u
m383 73033 5809 73013 VSS nch_18 l=0.65u w=1.3u
m384 73034 5809 73014 VSS nch_18 l=0.65u w=1.3u
m385 73035 5809 73015 VSS nch_18 l=0.65u w=1.3u
m386 73036 5809 73016 VSS nch_18 l=0.65u w=1.3u
m387 5800 5858 5786 VSS nch_18 l=0.55u w=0.65u
m388 73040 4994 73028 VSS nch_18 l=0.65u w=1.3u
m389 73041 4994 73029 VSS nch_18 l=0.65u w=1.3u
m390 73042 4994 73030 VSS nch_18 l=0.65u w=1.3u
m391 73043 4994 73031 VSS nch_18 l=0.65u w=1.3u
m392 5809 5823 5828 VSS nch_18 l=0.55u w=0.65u
m393 VSS 5809 73033 VSS nch_18 l=0.65u w=1.3u
m394 VSS 5809 73034 VSS nch_18 l=0.65u w=1.3u
m395 VSS 5809 73035 VSS nch_18 l=0.65u w=1.3u
m396 VSS 5809 73036 VSS nch_18 l=0.65u w=1.3u
m397 5786 5858 5800 VSS nch_18 l=0.55u w=0.65u
m398 5800 4994 73040 VSS nch_18 l=0.65u w=1.3u
m399 5800 4994 73041 VSS nch_18 l=0.65u w=1.3u
m400 5800 4994 73042 VSS nch_18 l=0.65u w=1.3u
m401 5800 4994 73043 VSS nch_18 l=0.65u w=1.3u
m402 73122 5809 5852 VSS nch_18 l=0.65u w=1.3u
m403 73123 5809 5852 VSS nch_18 l=0.65u w=1.3u
m404 73124 5809 5852 VSS nch_18 l=0.65u w=1.3u
m405 73125 5809 5852 VSS nch_18 l=0.65u w=1.3u
m406 5852 5823 5854 VSS nch_18 l=0.55u w=0.65u
m407 73133 5858 VSS VSS nch_18 l=0.65u w=1.3u
m408 73134 5858 VSS VSS nch_18 l=0.65u w=1.3u
m409 73135 5858 5858 VSS nch_18 l=0.65u w=1.3u
m410 73136 5858 5858 VSS nch_18 l=0.65u w=1.3u
m411 5854 5823 5852 VSS nch_18 l=0.55u w=0.65u
m412 73143 5809 73122 VSS nch_18 l=0.65u w=1.3u
m413 73144 5809 73123 VSS nch_18 l=0.65u w=1.3u
m414 73145 5809 73124 VSS nch_18 l=0.65u w=1.3u
m415 73146 5809 73125 VSS nch_18 l=0.65u w=1.3u
m416 73155 5858 73133 VSS nch_18 l=0.65u w=1.3u
m417 73156 5858 73134 VSS nch_18 l=0.65u w=1.3u
m418 73157 5858 73135 VSS nch_18 l=0.65u w=1.3u
m419 73158 5858 73136 VSS nch_18 l=0.65u w=1.3u
m420 5852 5823 5854 VSS nch_18 l=0.55u w=0.65u
m421 73162 5809 73143 VSS nch_18 l=0.65u w=1.3u
m422 73163 5809 73144 VSS nch_18 l=0.65u w=1.3u
m423 73164 5809 73145 VSS nch_18 l=0.65u w=1.3u
m424 73165 5809 73146 VSS nch_18 l=0.65u w=1.3u
m425 73173 5858 73155 VSS nch_18 l=0.65u w=1.3u
m426 73174 5858 73156 VSS nch_18 l=0.65u w=1.3u
m427 73175 5858 73157 VSS nch_18 l=0.65u w=1.3u
m428 73176 5858 73158 VSS nch_18 l=0.65u w=1.3u
m429 5854 5823 5852 VSS nch_18 l=0.55u w=0.65u
m430 VSS 5809 73162 VSS nch_18 l=0.65u w=1.3u
m431 VSS 5809 73163 VSS nch_18 l=0.65u w=1.3u
m432 VSS 5809 73164 VSS nch_18 l=0.65u w=1.3u
m433 VSS 5809 73165 VSS nch_18 l=0.65u w=1.3u
m434 5882 5858 73173 VSS nch_18 l=0.65u w=1.3u
m435 5882 5858 73174 VSS nch_18 l=0.65u w=1.3u
m436 5882 5858 73175 VSS nch_18 l=0.65u w=1.3u
m437 5882 5858 73176 VSS nch_18 l=0.65u w=1.3u
m438 6 PD VSS VSS nch l=0.04u w=0.4u
m439 VSS 6 8 VSS nch l=0.04u w=0.8u
m440 8 6 VSS VSS nch l=0.04u w=0.8u
m441 9 FREF 8 VSS nch l=0.04u w=0.62u
m442 10 FREF VSS VSS nch l=0.04u w=0.4u
m443 11 9 VSS VSS nch l=0.04u w=0.4u
m444 12 10 VSS VSS nch l=0.04u w=0.4u
m445 VSS 9 11 VSS nch l=0.04u w=0.4u
m446 VSS 10 12 VSS nch l=0.04u w=0.4u
m447 11 9 VSS VSS nch l=0.04u w=0.4u
m448 12 10 VSS VSS nch l=0.04u w=0.4u
m449 VSS 9 11 VSS nch l=0.04u w=0.4u
m450 VSS 10 12 VSS nch l=0.04u w=0.4u
m451 15 REFDIV[3] VSS VSS nch l=0.04u w=0.4u
m452 VSS 212 13 VSS nch l=0.04u w=0.8u
m453 VSS 30 14 VSS nch l=0.04u w=0.4u
m454 69143 110 VSS VSS nch l=0.04u w=0.8u
m455 69144 66 VSS VSS nch l=0.04u w=0.8u
m456 VSS REFDIV[4] 15 VSS nch l=0.04u w=0.4u
m457 13 212 VSS VSS nch l=0.04u w=0.8u
m458 17 91 69143 VSS nch l=0.04u w=0.8u
m459 18 94 69144 VSS nch l=0.04u w=0.8u
m460 15 REFDIV[5] VSS VSS nch l=0.04u w=0.4u
m461 16 11 13 VSS nch l=0.04u w=0.8u
m462 VSS 19 19 VSS nch l=0.04u w=0.8u
m463 69154 138 VSS VSS nch l=0.04u w=0.8u
m464 69155 77 21 VSS nch l=0.04u w=0.8u
m465 69156 130 VSS VSS nch l=0.04u w=0.8u
m466 69157 139 VSS VSS nch l=0.04u w=0.8u
m467 69158 78 22 VSS nch l=0.04u w=0.8u
m468 69159 140 VSS VSS nch l=0.04u w=0.8u
m469 69160 2616 VSS VSS nch l=0.04u w=0.8u
m470 69161 2616 VSS VSS nch l=0.04u w=0.8u
m471 VSS 23 23 VSS nch l=0.04u w=0.8u
m472 69162 141 VSS VSS nch l=0.04u w=0.8u
m473 69163 79 25 VSS nch l=0.04u w=0.8u
m474 69164 FRAC[0] VSS VSS nch l=0.04u w=0.8u
m475 43 60 VSS VSS nch l=0.04u w=0.4u
m476 44 61 VSS VSS nch l=0.04u w=0.4u
m477 VSS 109 26 VSS nch l=0.04u w=0.4u
m478 69165 81 27 VSS nch l=0.04u w=0.8u
m479 69166 132 VSS VSS nch l=0.04u w=0.8u
m480 46 4328 VSS VSS nch l=0.04u w=0.4u
m481 47 4328 VSS VSS nch l=0.04u w=0.4u
m482 69167 145 VSS VSS nch l=0.04u w=0.8u
m483 69168 82 28 VSS nch l=0.04u w=0.8u
m484 69169 146 VSS VSS nch l=0.04u w=0.8u
m485 69170 26 VSS VSS nch l=0.04u w=0.8u
m486 51 4328 VSS VSS nch l=0.04u w=0.4u
m487 52 4328 VSS VSS nch l=0.04u w=0.4u
m488 69171 141 VSS VSS nch l=0.04u w=0.8u
m489 69172 83 29 VSS nch l=0.04u w=0.8u
m490 69173 FRAC[0] VSS VSS nch l=0.04u w=0.8u
m491 69174 26 VSS VSS nch l=0.04u w=0.8u
m492 69175 84 30 VSS nch l=0.04u w=0.8u
m493 VSS 31 31 VSS nch l=0.04u w=0.8u
m494 VSS 34 34 VSS nch l=0.04u w=0.8u
m495 35 125 69154 VSS nch l=0.04u w=0.8u
m496 VSS 246 69155 VSS nch l=0.04u w=0.8u
m497 36 126 69156 VSS nch l=0.04u w=0.8u
m498 37 127 69157 VSS nch l=0.04u w=0.8u
m499 VSS 247 69158 VSS nch l=0.04u w=0.8u
m500 38 128 69159 VSS nch l=0.04u w=0.8u
m501 39 298 69160 VSS nch l=0.04u w=0.8u
m502 40 299 69161 VSS nch l=0.04u w=0.8u
m503 41 129 69162 VSS nch l=0.04u w=0.8u
m504 VSS 248 69163 VSS nch l=0.04u w=0.8u
m505 42 130 69164 VSS nch l=0.04u w=0.8u
m506 58 69 43 VSS nch l=0.04u w=0.4u
m507 59 70 44 VSS nch l=0.04u w=0.4u
m508 VSS 249 69165 VSS nch l=0.04u w=0.8u
m509 45 131 69166 VSS nch l=0.04u w=0.8u
m510 48 132 69167 VSS nch l=0.04u w=0.8u
m511 VSS 250 69168 VSS nch l=0.04u w=0.8u
m512 49 133 69169 VSS nch l=0.04u w=0.8u
m513 50 134 69170 VSS nch l=0.04u w=0.8u
m514 53 135 69171 VSS nch l=0.04u w=0.8u
m515 VSS 251 69172 VSS nch l=0.04u w=0.8u
m516 54 136 69173 VSS nch l=0.04u w=0.8u
m517 55 FBDIV[0] 69174 VSS nch l=0.04u w=0.8u
m518 VSS 2648 69175 VSS nch l=0.04u w=0.8u
m519 VSS 56 56 VSS nch l=0.04u w=0.8u
m520 VSS 20 VSS VSS nch l=0.26u w=0.8u
m521 VSS 24 VSS VSS nch l=0.26u w=0.8u
m522 67 91 VSS VSS nch l=0.04u w=0.4u
m523 68 94 VSS VSS nch l=0.04u w=0.4u
m524 69 43 58 VSS nch l=0.04u w=0.4u
m525 70 44 59 VSS nch l=0.04u w=0.4u
m526 75 REFDIV[1] VSS VSS nch l=0.04u w=0.4u
m527 76 16 VSS VSS nch l=0.04u w=0.4u
m528 80 4328 VSS VSS nch l=0.04u w=0.4u
m529 71 46 62 VSS nch l=0.04u w=0.4u
m530 72 47 63 VSS nch l=0.04u w=0.4u
m531 73 51 64 VSS nch l=0.04u w=0.4u
m532 74 52 65 VSS nch l=0.04u w=0.4u
m533 VSS 110 66 VSS nch l=0.04u w=0.4u
m534 VSS 32 VSS VSS nch l=0.26u w=0.8u
m535 VSS 33 VSS VSS nch l=0.26u w=0.8u
m536 89 110 67 VSS nch l=0.04u w=0.4u
m537 90 66 68 VSS nch l=0.04u w=0.4u
m538 VSS REFDIV[2] 75 VSS nch l=0.04u w=0.4u
m539 VSS 16 76 VSS nch l=0.04u w=0.4u
m540 92 125 VSS VSS nch l=0.04u w=0.4u
m541 69184 1159 77 VSS nch l=0.04u w=0.8u
m542 93 126 VSS VSS nch l=0.04u w=0.4u
m543 95 127 VSS VSS nch l=0.04u w=0.4u
m544 69185 1162 78 VSS nch l=0.04u w=0.8u
m545 96 128 VSS VSS nch l=0.04u w=0.4u
m546 97 39 VSS VSS nch l=0.04u w=0.4u
m547 98 40 VSS VSS nch l=0.04u w=0.4u
m548 99 129 VSS VSS nch l=0.04u w=0.4u
m549 69186 1165 79 VSS nch l=0.04u w=0.8u
m550 100 130 VSS VSS nch l=0.04u w=0.4u
m551 69187 131 81 VSS nch l=0.04u w=0.8u
m552 101 131 VSS VSS nch l=0.04u w=0.4u
m553 69188 4328 71 VSS nch l=0.04u w=0.12u
m554 69189 4328 72 VSS nch l=0.04u w=0.12u
m555 102 132 VSS VSS nch l=0.04u w=0.4u
m556 69190 1169 82 VSS nch l=0.04u w=0.8u
m557 103 133 VSS VSS nch l=0.04u w=0.4u
m558 104 134 VSS VSS nch l=0.04u w=0.4u
m559 69191 4328 73 VSS nch l=0.04u w=0.12u
m560 69192 4328 74 VSS nch l=0.04u w=0.12u
m561 105 135 VSS VSS nch l=0.04u w=0.4u
m562 69193 1173 83 VSS nch l=0.04u w=0.8u
m563 106 136 VSS VSS nch l=0.04u w=0.4u
m564 107 FBDIV[0] VSS VSS nch l=0.04u w=0.4u
m565 VSS 154 84 VSS nch l=0.04u w=0.4u
m566 108 DSMPD VSS VSS nch l=0.04u w=0.4u
m567 VSS 57 VSS VSS nch l=0.26u w=0.8u
m568 VSS 86 86 VSS nch l=0.04u w=0.8u
m569 VSS 87 87 VSS nch l=0.04u w=0.8u
m570 VSS 20 VSS VSS nch l=0.26u w=0.8u
m571 VSS 24 VSS VSS nch l=0.26u w=0.8u
m572 110 67 89 VSS nch l=0.04u w=0.4u
m573 66 68 90 VSS nch l=0.04u w=0.4u
m574 76 16 VSS VSS nch l=0.04u w=0.4u
m575 111 138 92 VSS nch l=0.04u w=0.4u
m576 69194 311 69184 VSS nch l=0.04u w=0.8u
m577 112 130 93 VSS nch l=0.04u w=0.4u
m578 113 139 95 VSS nch l=0.04u w=0.4u
m579 69195 312 69185 VSS nch l=0.04u w=0.8u
m580 114 140 96 VSS nch l=0.04u w=0.4u
m581 115 141 99 VSS nch l=0.04u w=0.4u
m582 69196 314 69186 VSS nch l=0.04u w=0.8u
m583 116 FRAC[0] 100 VSS nch l=0.04u w=0.4u
m584 69197 316 69187 VSS nch l=0.04u w=0.8u
m585 118 132 101 VSS nch l=0.04u w=0.4u
m586 VSS 143 69188 VSS nch l=0.04u w=0.12u
m587 VSS 144 69189 VSS nch l=0.04u w=0.12u
m588 119 145 102 VSS nch l=0.04u w=0.4u
m589 69198 317 69190 VSS nch l=0.04u w=0.8u
m590 120 146 103 VSS nch l=0.04u w=0.4u
m591 121 26 104 VSS nch l=0.04u w=0.4u
m592 VSS 147 69191 VSS nch l=0.04u w=0.12u
m593 VSS 148 69192 VSS nch l=0.04u w=0.12u
m594 122 141 105 VSS nch l=0.04u w=0.4u
m595 69199 319 69193 VSS nch l=0.04u w=0.8u
m596 123 FRAC[0] 106 VSS nch l=0.04u w=0.4u
m597 124 26 107 VSS nch l=0.04u w=0.4u
m598 69200 14 VSS VSS nch l=0.04u w=0.12u
m599 117 80 109 VSS nch l=0.04u w=0.4u
m600 VSS 32 VSS VSS nch l=0.26u w=0.8u
m601 VSS 33 VSS VSS nch l=0.26u w=0.8u
m602 VSS 16 76 VSS nch l=0.04u w=0.4u
m603 138 92 111 VSS nch l=0.04u w=0.4u
m604 VSS 160 69194 VSS nch l=0.04u w=0.8u
m605 130 93 112 VSS nch l=0.04u w=0.4u
m606 139 95 113 VSS nch l=0.04u w=0.4u
m607 VSS 162 69195 VSS nch l=0.04u w=0.8u
m608 140 96 114 VSS nch l=0.04u w=0.4u
m609 141 99 115 VSS nch l=0.04u w=0.4u
m610 VSS 163 69196 VSS nch l=0.04u w=0.8u
m611 FRAC[0] 100 116 VSS nch l=0.04u w=0.4u
m612 VSS 164 69197 VSS nch l=0.04u w=0.8u
m613 132 101 118 VSS nch l=0.04u w=0.4u
m614 143 71 VSS VSS nch l=0.04u w=0.4u
m615 144 72 VSS VSS nch l=0.04u w=0.4u
m616 145 102 119 VSS nch l=0.04u w=0.4u
m617 VSS 165 69198 VSS nch l=0.04u w=0.8u
m618 146 103 120 VSS nch l=0.04u w=0.4u
m619 26 104 121 VSS nch l=0.04u w=0.4u
m620 147 73 VSS VSS nch l=0.04u w=0.4u
m621 148 74 VSS VSS nch l=0.04u w=0.4u
m622 141 105 122 VSS nch l=0.04u w=0.4u
m623 VSS 166 69199 VSS nch l=0.04u w=0.8u
m624 FRAC[0] 106 123 VSS nch l=0.04u w=0.4u
m625 26 107 124 VSS nch l=0.04u w=0.4u
m626 69201 75 VSS VSS nch l=0.04u w=0.8u
m627 154 270 69200 VSS nch l=0.04u w=0.12u
m628 150 4328 VSS VSS nch l=0.04u w=0.4u
m629 151 4328 VSS VSS nch l=0.04u w=0.4u
m630 152 4328 VSS VSS nch l=0.04u w=0.4u
m631 153 4328 VSS VSS nch l=0.04u w=0.4u
m632 69202 4328 117 VSS nch l=0.04u w=0.12u
m633 69203 14 VSS VSS nch l=0.04u w=0.8u
m634 VSS 57 VSS VSS nch l=0.26u w=0.8u
m635 VSS 85 VSS VSS nch l=0.26u w=0.8u
m636 VSS 88 VSS VSS nch l=0.26u w=0.8u
m637 VSS 20 VSS VSS nch l=0.26u w=0.8u
m638 VSS 24 VSS VSS nch l=0.26u w=0.8u
m639 156 4328 VSS VSS nch l=0.04u w=0.4u
m640 157 4328 VSS VSS nch l=0.04u w=0.4u
m641 76 16 VSS VSS nch l=0.04u w=0.4u
m642 149 15 69201 VSS nch l=0.04u w=0.8u
m643 158 886 154 VSS nch l=0.04u w=0.4u
m644 VSS 177 69202 VSS nch l=0.04u w=0.12u
m645 155 108 69203 VSS nch l=0.04u w=0.8u
m646 VSS 32 VSS VSS nch l=0.26u w=0.8u
m647 VSS 33 VSS VSS nch l=0.26u w=0.8u
m648 VSS 16 76 VSS nch l=0.04u w=0.4u
m649 VSS 57 VSS VSS nch l=0.26u w=0.8u
m650 69219 89 159 VSS nch l=0.04u w=0.8u
m651 VSS 194 160 VSS nch l=0.04u w=0.4u
m652 69220 90 161 VSS nch l=0.04u w=0.8u
m653 VSS 195 162 VSS nch l=0.04u w=0.4u
m654 VSS 196 163 VSS nch l=0.04u w=0.4u
m655 177 117 VSS VSS nch l=0.04u w=0.4u
m656 VSS 197 164 VSS nch l=0.04u w=0.4u
m657 169 4328 143 VSS nch l=0.04u w=0.4u
m658 170 4328 144 VSS nch l=0.04u w=0.4u
m659 VSS 198 165 VSS nch l=0.04u w=0.4u
m660 171 4328 147 VSS nch l=0.04u w=0.4u
m661 172 4328 148 VSS nch l=0.04u w=0.4u
m662 VSS 199 166 VSS nch l=0.04u w=0.4u
m663 173 150 167 VSS nch l=0.04u w=0.4u
m664 174 151 168 VSS nch l=0.04u w=0.4u
m665 175 152 97 VSS nch l=0.04u w=0.4u
m666 176 153 98 VSS nch l=0.04u w=0.4u
m667 VSS 85 VSS VSS nch l=0.26u w=0.8u
m668 VSS 88 VSS VSS nch l=0.26u w=0.8u
m669 VSS 20 VSS VSS nch l=0.26u w=0.8u
m670 VSS 24 VSS VSS nch l=0.26u w=0.8u
m671 76 16 VSS VSS nch l=0.04u w=0.4u
m672 191 156 58 VSS nch l=0.04u w=0.4u
m673 192 157 59 VSS nch l=0.04u w=0.4u
m674 VSS 110 69219 VSS nch l=0.04u w=0.8u
m675 VSS 293 69220 VSS nch l=0.04u w=0.8u
m676 69221 46 169 VSS nch l=0.04u w=0.12u
m677 69222 47 170 VSS nch l=0.04u w=0.12u
m678 69223 51 171 VSS nch l=0.04u w=0.12u
m679 69224 52 172 VSS nch l=0.04u w=0.12u
m680 193 149 VSS VSS nch l=0.04u w=0.4u
m681 69225 217 158 VSS nch l=0.04u w=0.8u
m682 69226 4328 173 VSS nch l=0.04u w=0.12u
m683 69227 4328 174 VSS nch l=0.04u w=0.12u
m684 69228 111 178 VSS nch l=0.04u w=0.8u
m685 69229 112 179 VSS nch l=0.04u w=0.8u
m686 69230 113 180 VSS nch l=0.04u w=0.8u
m687 69231 114 181 VSS nch l=0.04u w=0.8u
m688 69232 4328 175 VSS nch l=0.04u w=0.12u
m689 69233 4328 176 VSS nch l=0.04u w=0.12u
m690 69234 115 182 VSS nch l=0.04u w=0.8u
m691 69235 116 183 VSS nch l=0.04u w=0.8u
m692 69236 118 184 VSS nch l=0.04u w=0.8u
m693 69237 119 185 VSS nch l=0.04u w=0.8u
m694 69238 120 186 VSS nch l=0.04u w=0.8u
m695 69239 121 187 VSS nch l=0.04u w=0.8u
m696 69240 122 188 VSS nch l=0.04u w=0.8u
m697 69241 123 189 VSS nch l=0.04u w=0.8u
m698 69242 124 190 VSS nch l=0.04u w=0.8u
m699 200 155 VSS VSS nch l=0.04u w=0.4u
m700 VSS 32 VSS VSS nch l=0.26u w=0.8u
m701 VSS 33 VSS VSS nch l=0.26u w=0.8u
m702 VSS 16 76 VSS nch l=0.04u w=0.4u
m703 VSS 57 VSS VSS nch l=0.26u w=0.8u
m704 69243 4328 191 VSS nch l=0.04u w=0.12u
m705 69244 4328 192 VSS nch l=0.04u w=0.12u
m706 VSS 202 69221 VSS nch l=0.04u w=0.12u
m707 VSS 203 69222 VSS nch l=0.04u w=0.12u
m708 VSS 204 69223 VSS nch l=0.04u w=0.12u
m709 VSS 205 69224 VSS nch l=0.04u w=0.12u
m710 VSS 2648 69225 VSS nch l=0.04u w=0.8u
m711 VSS 207 69226 VSS nch l=0.04u w=0.12u
m712 VSS 208 69227 VSS nch l=0.04u w=0.12u
m713 VSS 21 69228 VSS nch l=0.04u w=0.8u
m714 69245 610 194 VSS nch l=0.04u w=0.8u
m715 VSS 110 69229 VSS nch l=0.04u w=0.8u
m716 VSS 22 69230 VSS nch l=0.04u w=0.8u
m717 69246 611 195 VSS nch l=0.04u w=0.8u
m718 VSS 313 69231 VSS nch l=0.04u w=0.8u
m719 VSS 210 69232 VSS nch l=0.04u w=0.12u
m720 VSS 211 69233 VSS nch l=0.04u w=0.12u
m721 VSS 25 69234 VSS nch l=0.04u w=0.8u
m722 69247 612 196 VSS nch l=0.04u w=0.8u
m723 VSS 315 69235 VSS nch l=0.04u w=0.8u
m724 201 4328 177 VSS nch l=0.04u w=0.4u
m725 69248 613 197 VSS nch l=0.04u w=0.8u
m726 VSS 27 69236 VSS nch l=0.04u w=0.8u
m727 VSS 28 69237 VSS nch l=0.04u w=0.8u
m728 69249 614 198 VSS nch l=0.04u w=0.8u
m729 VSS 131 69238 VSS nch l=0.04u w=0.8u
m730 VSS 318 69239 VSS nch l=0.04u w=0.8u
m731 VSS 29 69240 VSS nch l=0.04u w=0.8u
m732 69250 615 199 VSS nch l=0.04u w=0.8u
m733 VSS 131 69241 VSS nch l=0.04u w=0.8u
m734 VSS 318 69242 VSS nch l=0.04u w=0.8u
m735 VSS 85 VSS VSS nch l=0.26u w=0.8u
m736 VSS 88 VSS VSS nch l=0.26u w=0.8u
m737 VSS 20 VSS VSS nch l=0.26u w=0.8u
m738 VSS 24 VSS VSS nch l=0.26u w=0.8u
m739 VSS 214 69243 VSS nch l=0.04u w=0.12u
m740 VSS 215 69244 VSS nch l=0.04u w=0.12u
m741 202 169 VSS VSS nch l=0.04u w=0.4u
m742 203 170 VSS VSS nch l=0.04u w=0.4u
m743 204 171 VSS VSS nch l=0.04u w=0.4u
m744 205 172 VSS VSS nch l=0.04u w=0.4u
m745 69251 158 VSS VSS nch l=0.04u w=0.24u
m746 69252 159 VSS VSS nch l=0.04u w=0.8u
m747 207 173 VSS VSS nch l=0.04u w=0.4u
m748 208 174 VSS VSS nch l=0.04u w=0.4u
m749 69253 903 69245 VSS nch l=0.04u w=0.8u
m750 69254 161 VSS VSS nch l=0.04u w=0.8u
m751 69255 904 69246 VSS nch l=0.04u w=0.8u
m752 210 175 VSS VSS nch l=0.04u w=0.4u
m753 211 176 VSS VSS nch l=0.04u w=0.4u
m754 69256 905 69247 VSS nch l=0.04u w=0.8u
m755 69257 80 201 VSS nch l=0.04u w=0.12u
m756 69258 906 69248 VSS nch l=0.04u w=0.8u
m757 69259 907 69249 VSS nch l=0.04u w=0.8u
m758 69260 908 69250 VSS nch l=0.04u w=0.8u
m759 212 PD VSS VSS nch l=0.04u w=0.4u
m760 VSS 32 VSS VSS nch l=0.26u w=0.8u
m761 VSS 33 VSS VSS nch l=0.26u w=0.8u
m762 69261 155 VSS VSS nch l=0.04u w=0.8u
m763 VSS 57 VSS VSS nch l=0.26u w=0.8u
m764 214 191 VSS VSS nch l=0.04u w=0.4u
m765 215 192 VSS VSS nch l=0.04u w=0.4u
m766 216 236 VSS VSS nch l=0.04u w=0.4u
m767 217 886 69251 VSS nch l=0.04u w=0.24u
m768 206 17 69252 VSS nch l=0.04u w=0.8u
m769 VSS 1190 69253 VSS nch l=0.04u w=0.8u
m770 209 18 69254 VSS nch l=0.04u w=0.8u
m771 VSS 1191 69255 VSS nch l=0.04u w=0.8u
m772 VSS 1192 69256 VSS nch l=0.04u w=0.8u
m773 VSS 241 69257 VSS nch l=0.04u w=0.12u
m774 VSS 1193 69258 VSS nch l=0.04u w=0.8u
m775 VSS 1194 69259 VSS nch l=0.04u w=0.8u
m776 VSS 1195 69260 VSS nch l=0.04u w=0.8u
m777 VSS 193 212 VSS nch l=0.04u w=0.4u
m778 VSS 85 VSS VSS nch l=0.26u w=0.8u
m779 VSS 88 VSS VSS nch l=0.26u w=0.8u
m780 69262 178 VSS VSS nch l=0.04u w=0.8u
m781 69263 179 VSS VSS nch l=0.04u w=0.8u
m782 69264 180 VSS VSS nch l=0.04u w=0.8u
m783 69265 181 VSS VSS nch l=0.04u w=0.8u
m784 69266 182 VSS VSS nch l=0.04u w=0.8u
m785 69267 183 VSS VSS nch l=0.04u w=0.8u
m786 69268 184 VSS VSS nch l=0.04u w=0.8u
m787 69269 185 VSS VSS nch l=0.04u w=0.8u
m788 69270 186 VSS VSS nch l=0.04u w=0.8u
m789 69271 187 VSS VSS nch l=0.04u w=0.8u
m790 69272 188 VSS VSS nch l=0.04u w=0.8u
m791 69273 189 VSS VSS nch l=0.04u w=0.8u
m792 69274 190 VSS VSS nch l=0.04u w=0.8u
m793 231 232 VSS VSS nch l=0.04u w=0.8u
m794 234 233 VSS VSS nch l=0.04u w=0.8u
m795 213 FBDIV[0] 69261 VSS nch l=0.04u w=0.8u
m796 VSS 20 VSS VSS nch l=0.26u w=0.8u
m797 VSS 24 VSS VSS nch l=0.26u w=0.8u
m798 VDDREF 270 217 VSS nch l=0.04u w=0.4u
m799 241 201 VSS VSS nch l=0.04u w=0.4u
m800 242 4328 VSS VSS nch l=0.04u w=0.4u
m801 243 4328 VSS VSS nch l=0.04u w=0.4u
m802 244 4328 VSS VSS nch l=0.04u w=0.4u
m803 245 4328 VSS VSS nch l=0.04u w=0.4u
m804 237 4328 207 VSS nch l=0.04u w=0.4u
m805 238 4328 208 VSS nch l=0.04u w=0.4u
m806 218 35 69262 VSS nch l=0.04u w=0.8u
m807 219 36 69263 VSS nch l=0.04u w=0.8u
m808 220 37 69264 VSS nch l=0.04u w=0.8u
m809 221 38 69265 VSS nch l=0.04u w=0.8u
m810 239 4328 210 VSS nch l=0.04u w=0.4u
m811 240 4328 211 VSS nch l=0.04u w=0.4u
m812 222 41 69266 VSS nch l=0.04u w=0.8u
m813 223 42 69267 VSS nch l=0.04u w=0.8u
m814 224 45 69268 VSS nch l=0.04u w=0.8u
m815 225 48 69269 VSS nch l=0.04u w=0.8u
m816 226 49 69270 VSS nch l=0.04u w=0.8u
m817 227 50 69271 VSS nch l=0.04u w=0.8u
m818 228 53 69272 VSS nch l=0.04u w=0.8u
m819 229 54 69273 VSS nch l=0.04u w=0.8u
m820 230 55 69274 VSS nch l=0.04u w=0.8u
m821 VSS 57 VSS VSS nch l=0.26u w=0.8u
m822 257 4328 214 VSS nch l=0.04u w=0.4u
m823 258 4328 215 VSS nch l=0.04u w=0.4u
m824 235 259 236 VSS nch l=0.04u w=0.4u
m825 VSS 85 VSS VSS nch l=0.26u w=0.8u
m826 VSS 88 VSS VSS nch l=0.26u w=0.8u
m827 260 89 VSS VSS nch l=0.04u w=0.4u
m828 69275 150 237 VSS nch l=0.04u w=0.12u
m829 69276 151 238 VSS nch l=0.04u w=0.12u
m830 VSS 353 246 VSS nch l=0.04u w=0.4u
m831 261 90 VSS VSS nch l=0.04u w=0.4u
m832 VSS 356 247 VSS nch l=0.04u w=0.4u
m833 69277 152 239 VSS nch l=0.04u w=0.12u
m834 69278 153 240 VSS nch l=0.04u w=0.12u
m835 VSS 361 248 VSS nch l=0.04u w=0.4u
m836 VSS 363 249 VSS nch l=0.04u w=0.4u
m837 VSS 366 250 VSS nch l=0.04u w=0.4u
m838 VSS 370 251 VSS nch l=0.04u w=0.4u
m839 236 212 VSS VSS nch l=0.04u w=0.4u
m840 VSS 20 VSS VSS nch l=0.26u w=0.8u
m841 VSS 24 VSS VSS nch l=0.26u w=0.8u
m842 VSS 252 252 VSS nch l=0.04u w=0.8u
m843 VSS 255 255 VSS nch l=0.04u w=0.8u
m844 69280 200 VSS VSS nch l=0.04u w=0.8u
m845 69282 156 257 VSS nch l=0.04u w=0.12u
m846 69283 157 258 VSS nch l=0.04u w=0.12u
m847 259 236 235 VSS nch l=0.04u w=0.4u
m848 270 886 VSS VSS nch l=0.04u w=0.4u
m849 271 110 260 VSS nch l=0.04u w=0.4u
m850 VSS 292 69275 VSS nch l=0.04u w=0.12u
m851 VSS 126 69276 VSS nch l=0.04u w=0.12u
m852 272 293 261 VSS nch l=0.04u w=0.4u
m853 VSS 294 69277 VSS nch l=0.04u w=0.12u
m854 VSS 130 69278 VSS nch l=0.04u w=0.12u
m855 266 242 262 VSS nch l=0.04u w=0.4u
m856 267 243 263 VSS nch l=0.04u w=0.4u
m857 268 244 264 VSS nch l=0.04u w=0.4u
m858 269 245 134 VSS nch l=0.04u w=0.4u
m859 273 111 VSS VSS nch l=0.04u w=0.4u
m860 275 112 VSS VSS nch l=0.04u w=0.4u
m861 276 113 VSS VSS nch l=0.04u w=0.4u
m862 278 114 VSS VSS nch l=0.04u w=0.4u
m863 279 115 VSS VSS nch l=0.04u w=0.4u
m864 281 116 VSS VSS nch l=0.04u w=0.4u
m865 283 118 VSS VSS nch l=0.04u w=0.4u
m866 284 119 VSS VSS nch l=0.04u w=0.4u
m867 286 120 VSS VSS nch l=0.04u w=0.4u
m868 287 121 VSS VSS nch l=0.04u w=0.4u
m869 288 122 VSS VSS nch l=0.04u w=0.4u
m870 290 123 VSS VSS nch l=0.04u w=0.4u
m871 291 124 VSS VSS nch l=0.04u w=0.4u
m872 265 241 69280 VSS nch l=0.04u w=0.8u
m873 VSS 57 VSS VSS nch l=0.26u w=0.8u
m874 VSS 85 VSS VSS nch l=0.26u w=0.8u
m875 VSS 88 VSS VSS nch l=0.26u w=0.8u
m876 VSS 304 69282 VSS nch l=0.04u w=0.12u
m877 VSS 305 69283 VSS nch l=0.04u w=0.12u
m878 110 260 271 VSS nch l=0.04u w=0.4u
m879 292 237 VSS VSS nch l=0.04u w=0.4u
m880 126 238 VSS VSS nch l=0.04u w=0.4u
m881 VSS 20 VSS VSS nch l=0.26u w=0.8u
m882 293 261 272 VSS nch l=0.04u w=0.4u
m883 294 239 VSS VSS nch l=0.04u w=0.4u
m884 130 240 VSS VSS nch l=0.04u w=0.4u
m885 VSS 24 VSS VSS nch l=0.26u w=0.8u
m886 69292 4328 266 VSS nch l=0.04u w=0.12u
m887 69293 4328 267 VSS nch l=0.04u w=0.12u
m888 69294 4328 268 VSS nch l=0.04u w=0.12u
m889 69295 4328 269 VSS nch l=0.04u w=0.12u
m890 VSS 253 VSS VSS nch l=0.26u w=0.8u
m891 VSS 254 VSS VSS nch l=0.26u w=0.8u
m892 296 21 273 VSS nch l=0.04u w=0.4u
m893 168 110 275 VSS nch l=0.04u w=0.4u
m894 297 22 276 VSS nch l=0.04u w=0.4u
m895 299 313 278 VSS nch l=0.04u w=0.4u
m896 127 25 279 VSS nch l=0.04u w=0.4u
m897 128 315 281 VSS nch l=0.04u w=0.4u
m898 109 27 283 VSS nch l=0.04u w=0.4u
m899 263 28 284 VSS nch l=0.04u w=0.4u
m900 302 131 286 VSS nch l=0.04u w=0.4u
m901 145 318 287 VSS nch l=0.04u w=0.4u
m902 134 29 288 VSS nch l=0.04u w=0.4u
m903 146 131 290 VSS nch l=0.04u w=0.4u
m904 141 318 291 VSS nch l=0.04u w=0.4u
m905 303 485 VSS VSS nch l=0.04u w=0.4u
m906 304 257 VSS VSS nch l=0.04u w=0.4u
m907 305 258 VSS VSS nch l=0.04u w=0.4u
m908 306 377 VSS VSS nch l=0.04u w=0.4u
m909 307 308 VSS VSS nch l=0.04u w=0.8u
m910 309 310 VSS VSS nch l=0.04u w=0.8u
m911 VSS 323 69292 VSS nch l=0.04u w=0.12u
m912 VSS 324 69293 VSS nch l=0.04u w=0.12u
m913 VSS 325 69294 VSS nch l=0.04u w=0.12u
m914 VSS 326 69295 VSS nch l=0.04u w=0.12u
m915 VSS 327 LOCK VSS nch l=0.04u w=0.4u
m916 21 273 296 VSS nch l=0.04u w=0.4u
m917 110 275 168 VSS nch l=0.04u w=0.4u
m918 22 276 297 VSS nch l=0.04u w=0.4u
m919 313 278 299 VSS nch l=0.04u w=0.4u
m920 25 279 127 VSS nch l=0.04u w=0.4u
m921 315 281 128 VSS nch l=0.04u w=0.4u
m922 27 283 109 VSS nch l=0.04u w=0.4u
m923 28 284 263 VSS nch l=0.04u w=0.4u
m924 131 286 302 VSS nch l=0.04u w=0.4u
m925 318 287 145 VSS nch l=0.04u w=0.4u
m926 29 288 134 VSS nch l=0.04u w=0.4u
m927 131 290 146 VSS nch l=0.04u w=0.4u
m928 318 291 141 VSS nch l=0.04u w=0.4u
m929 VSS 485 303 VSS nch l=0.04u w=0.4u
m930 167 328 274 VSS nch l=0.04u w=0.4u
m931 298 329 277 VSS nch l=0.04u w=0.4u
m932 300 330 280 VSS nch l=0.04u w=0.4u
m933 301 331 282 VSS nch l=0.04u w=0.4u
m934 63 332 285 VSS nch l=0.04u w=0.4u
m935 65 333 289 VSS nch l=0.04u w=0.4u
m936 69297 265 VSS VSS nch l=0.04u w=0.8u
m937 VSS 57 VSS VSS nch l=0.26u w=0.8u
m938 VSS 85 VSS VSS nch l=0.26u w=0.8u
m939 VSS 88 VSS VSS nch l=0.26u w=0.8u
m940 VSS 253 VSS VSS nch l=0.26u w=0.8u
m941 VSS 254 VSS VSS nch l=0.26u w=0.8u
m942 323 266 VSS VSS nch l=0.04u w=0.4u
m943 324 267 VSS VSS nch l=0.04u w=0.4u
m944 325 268 VSS VSS nch l=0.04u w=0.4u
m945 326 269 VSS VSS nch l=0.04u w=0.4u
m946 303 485 VSS VSS nch l=0.04u w=0.4u
m947 328 274 167 VSS nch l=0.04u w=0.4u
m948 329 277 298 VSS nch l=0.04u w=0.4u
m949 330 280 300 VSS nch l=0.04u w=0.4u
m950 331 282 301 VSS nch l=0.04u w=0.4u
m951 332 285 63 VSS nch l=0.04u w=0.4u
m952 333 289 65 VSS nch l=0.04u w=0.4u
m953 320 213 69297 VSS nch l=0.04u w=0.8u
m954 334 335 VSS VSS nch l=0.04u w=0.8u
m955 VSS 304 321 VSS nch l=0.04u w=0.4u
m956 VSS 305 322 VSS nch l=0.04u w=0.4u
m957 69322 377 VSS VSS nch l=0.04u w=0.8u
m958 VSS 485 303 VSS nch l=0.04u w=0.4u
m959 69325 378 327 VSS nch l=0.04u w=0.8u
m960 69326 415 VSS VSS nch l=0.04u w=0.8u
m961 VSS 311 328 VSS nch l=0.04u w=0.4u
m962 69327 379 VSS VSS nch l=0.04u w=0.8u
m963 VSS 312 329 VSS nch l=0.04u w=0.4u
m964 VSS 314 330 VSS nch l=0.04u w=0.4u
m965 VSS 316 331 VSS nch l=0.04u w=0.4u
m966 VSS 317 332 VSS nch l=0.04u w=0.4u
m967 VSS 319 333 VSS nch l=0.04u w=0.4u
m968 VSS 85 VSS VSS nch l=0.26u w=0.8u
m969 VSS 88 VSS VSS nch l=0.26u w=0.8u
m970 VSS 253 VSS VSS nch l=0.26u w=0.8u
m971 VSS 254 VSS VSS nch l=0.26u w=0.8u
m972 346 321 VSS VSS nch l=0.04u w=0.4u
m973 347 322 VSS VSS nch l=0.04u w=0.4u
m974 336 REFDIV[0] 69322 VSS nch l=0.04u w=0.8u
m975 348 4328 323 VSS nch l=0.04u w=0.4u
m976 349 4328 324 VSS nch l=0.04u w=0.4u
m977 350 4328 325 VSS nch l=0.04u w=0.4u
m978 351 4328 326 VSS nch l=0.04u w=0.4u
m979 VSS 2648 69325 VSS nch l=0.04u w=0.8u
m980 337 395 69326 VSS nch l=0.04u w=0.8u
m981 338 398 69327 VSS nch l=0.04u w=0.8u
m982 VSS 339 339 VSS nch l=0.04u w=0.8u
m983 69329 458 VSS VSS nch l=0.04u w=0.8u
m984 69330 442 VSS VSS nch l=0.04u w=0.8u
m985 69331 139 VSS VSS nch l=0.04u w=0.8u
m986 69332 459 VSS VSS nch l=0.04u w=0.8u
m987 69333 2616 VSS VSS nch l=0.04u w=0.8u
m988 69334 2616 VSS VSS nch l=0.04u w=0.8u
m989 VSS 341 341 VSS nch l=0.04u w=0.8u
m990 69335 460 VSS VSS nch l=0.04u w=0.8u
m991 69336 FRAC[1] VSS VSS nch l=0.04u w=0.8u
m992 VSS 412 343 VSS nch l=0.04u w=0.4u
m993 69337 443 VSS VSS nch l=0.04u w=0.8u
m994 69338 462 VSS VSS nch l=0.04u w=0.8u
m995 69339 264 VSS VSS nch l=0.04u w=0.8u
m996 69340 343 VSS VSS nch l=0.04u w=0.8u
m997 69341 460 VSS VSS nch l=0.04u w=0.8u
m998 69342 FRAC[1] VSS VSS nch l=0.04u w=0.8u
m999 69343 343 VSS VSS nch l=0.04u w=0.8u
m1000 VSS 344 344 VSS nch l=0.04u w=0.8u
m1001 374 373 VSS VSS nch l=0.04u w=0.8u
m1002 375 376 VSS VSS nch l=0.04u w=0.8u
m1003 69345 242 348 VSS nch l=0.04u w=0.12u
m1004 69346 243 349 VSS nch l=0.04u w=0.12u
m1005 69347 244 350 VSS nch l=0.04u w=0.12u
m1006 69348 245 351 VSS nch l=0.04u w=0.12u
m1007 377 457 VSS VSS nch l=0.04u w=0.4u
m1008 352 437 69329 VSS nch l=0.04u w=0.8u
m1009 69349 530 353 VSS nch l=0.04u w=0.8u
m1010 354 438 69330 VSS nch l=0.04u w=0.8u
m1011 355 439 69331 VSS nch l=0.04u w=0.8u
m1012 69350 533 356 VSS nch l=0.04u w=0.8u
m1013 357 440 69332 VSS nch l=0.04u w=0.8u
m1014 358 597 69333 VSS nch l=0.04u w=0.8u
m1015 359 598 69334 VSS nch l=0.04u w=0.8u
m1016 360 441 69335 VSS nch l=0.04u w=0.8u
m1017 69351 536 361 VSS nch l=0.04u w=0.8u
m1018 362 442 69336 VSS nch l=0.04u w=0.8u
m1019 69352 538 363 VSS nch l=0.04u w=0.8u
m1020 364 131 69337 VSS nch l=0.04u w=0.8u
m1021 365 443 69338 VSS nch l=0.04u w=0.8u
m1022 69353 541 366 VSS nch l=0.04u w=0.8u
m1023 367 391 69339 VSS nch l=0.04u w=0.8u
m1024 368 444 69340 VSS nch l=0.04u w=0.8u
m1025 369 445 69341 VSS nch l=0.04u w=0.8u
m1026 69354 545 370 VSS nch l=0.04u w=0.8u
m1027 371 392 69342 VSS nch l=0.04u w=0.8u
m1028 372 FBDIV[1] 69343 VSS nch l=0.04u w=0.8u
m1029 VSS 253 VSS VSS nch l=0.26u w=0.8u
m1030 VSS 254 VSS VSS nch l=0.26u w=0.8u
m1031 385 4328 VSS VSS nch l=0.04u w=0.4u
m1032 386 4328 VSS VSS nch l=0.04u w=0.4u
m1033 VSS 391 69345 VSS nch l=0.04u w=0.12u
m1034 VSS 132 69346 VSS nch l=0.04u w=0.12u
m1035 VSS 392 69347 VSS nch l=0.04u w=0.12u
m1036 VSS 135 69348 VSS nch l=0.04u w=0.12u
m1037 69357 306 VSS VSS nch l=0.04u w=0.8u
m1038 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1039 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1040 VSS 457 377 VSS nch l=0.04u w=0.4u
m1041 VSS 416 378 VSS nch l=0.04u w=0.4u
m1042 388 395 VSS VSS nch l=0.04u w=0.4u
m1043 VSS 418 69349 VSS nch l=0.04u w=0.8u
m1044 389 398 VSS VSS nch l=0.04u w=0.4u
m1045 VSS 421 69350 VSS nch l=0.04u w=0.8u
m1046 VSS 424 69351 VSS nch l=0.04u w=0.8u
m1047 VSS 427 69352 VSS nch l=0.04u w=0.8u
m1048 VSS 430 69353 VSS nch l=0.04u w=0.8u
m1049 VSS 434 69354 VSS nch l=0.04u w=0.8u
m1050 390 4328 VSS VSS nch l=0.04u w=0.4u
m1051 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1052 VSS 1918 379 VSS nch l=0.04u w=0.4u
m1053 VSS 381 381 VSS nch l=0.04u w=0.8u
m1054 VSS 382 382 VSS nch l=0.04u w=0.8u
m1055 391 348 VSS VSS nch l=0.04u w=0.4u
m1056 132 349 VSS VSS nch l=0.04u w=0.4u
m1057 392 350 VSS VSS nch l=0.04u w=0.4u
m1058 135 351 VSS VSS nch l=0.04u w=0.4u
m1059 387 235 69357 VSS nch l=0.04u w=0.8u
m1060 377 457 VSS VSS nch l=0.04u w=0.4u
m1061 69359 LOCK VSS VSS nch l=0.04u w=0.12u
m1062 393 415 388 VSS nch l=0.04u w=0.4u
m1063 394 379 389 VSS nch l=0.04u w=0.4u
m1064 396 437 VSS VSS nch l=0.04u w=0.4u
m1065 397 438 VSS VSS nch l=0.04u w=0.4u
m1066 399 439 VSS VSS nch l=0.04u w=0.4u
m1067 400 440 VSS VSS nch l=0.04u w=0.4u
m1068 401 358 VSS VSS nch l=0.04u w=0.4u
m1069 402 359 VSS VSS nch l=0.04u w=0.4u
m1070 403 441 VSS VSS nch l=0.04u w=0.4u
m1071 404 442 VSS VSS nch l=0.04u w=0.4u
m1072 405 131 VSS VSS nch l=0.04u w=0.4u
m1073 406 443 VSS VSS nch l=0.04u w=0.4u
m1074 407 391 VSS VSS nch l=0.04u w=0.4u
m1075 408 444 VSS VSS nch l=0.04u w=0.4u
m1076 409 445 VSS VSS nch l=0.04u w=0.4u
m1077 410 392 VSS VSS nch l=0.04u w=0.4u
m1078 411 FBDIV[1] VSS VSS nch l=0.04u w=0.4u
m1079 VSS 253 VSS VSS nch l=0.26u w=0.8u
m1080 VSS 254 VSS VSS nch l=0.26u w=0.8u
m1081 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1082 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1083 413 385 304 VSS nch l=0.04u w=0.4u
m1084 414 386 305 VSS nch l=0.04u w=0.4u
m1085 VSS 457 377 VSS nch l=0.04u w=0.4u
m1086 416 561 69359 VSS nch l=0.04u w=0.12u
m1087 415 388 393 VSS nch l=0.04u w=0.4u
m1088 379 389 394 VSS nch l=0.04u w=0.4u
m1089 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1090 417 458 396 VSS nch l=0.04u w=0.4u
m1091 69360 274 VSS VSS nch l=0.04u w=0.8u
m1092 419 442 397 VSS nch l=0.04u w=0.4u
m1093 420 139 399 VSS nch l=0.04u w=0.4u
m1094 69361 277 VSS VSS nch l=0.04u w=0.8u
m1095 422 459 400 VSS nch l=0.04u w=0.4u
m1096 423 460 403 VSS nch l=0.04u w=0.4u
m1097 69362 280 VSS VSS nch l=0.04u w=0.8u
m1098 425 FRAC[1] 404 VSS nch l=0.04u w=0.4u
m1099 69363 282 VSS VSS nch l=0.04u w=0.8u
m1100 428 443 405 VSS nch l=0.04u w=0.4u
m1101 429 462 406 VSS nch l=0.04u w=0.4u
m1102 69364 285 VSS VSS nch l=0.04u w=0.8u
m1103 431 264 407 VSS nch l=0.04u w=0.4u
m1104 432 343 408 VSS nch l=0.04u w=0.4u
m1105 433 460 409 VSS nch l=0.04u w=0.4u
m1106 69365 289 VSS VSS nch l=0.04u w=0.8u
m1107 435 FRAC[1] 410 VSS nch l=0.04u w=0.4u
m1108 436 343 411 VSS nch l=0.04u w=0.4u
m1109 426 390 412 VSS nch l=0.04u w=0.4u
m1110 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1111 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1112 447 448 VSS VSS nch l=0.04u w=0.8u
m1113 450 449 VSS VSS nch l=0.04u w=0.8u
m1114 69367 4328 413 VSS nch l=0.04u w=0.12u
m1115 69368 4328 414 VSS nch l=0.04u w=0.12u
m1116 451 4328 VSS VSS nch l=0.04u w=0.4u
m1117 452 4328 VSS VSS nch l=0.04u w=0.4u
m1118 453 4328 VSS VSS nch l=0.04u w=0.4u
m1119 454 4328 VSS VSS nch l=0.04u w=0.4u
m1120 69369 387 VSS VSS nch l=0.04u w=0.8u
m1121 456 605 416 VSS nch l=0.04u w=0.4u
m1122 458 396 417 VSS nch l=0.04u w=0.4u
m1123 418 311 69360 VSS nch l=0.04u w=0.8u
m1124 442 397 419 VSS nch l=0.04u w=0.4u
m1125 139 399 420 VSS nch l=0.04u w=0.4u
m1126 421 312 69361 VSS nch l=0.04u w=0.8u
m1127 459 400 422 VSS nch l=0.04u w=0.4u
m1128 460 403 423 VSS nch l=0.04u w=0.4u
m1129 424 314 69362 VSS nch l=0.04u w=0.8u
m1130 FRAC[1] 404 425 VSS nch l=0.04u w=0.4u
m1131 427 316 69363 VSS nch l=0.04u w=0.8u
m1132 443 405 428 VSS nch l=0.04u w=0.4u
m1133 462 406 429 VSS nch l=0.04u w=0.4u
m1134 430 317 69364 VSS nch l=0.04u w=0.8u
m1135 264 407 431 VSS nch l=0.04u w=0.4u
m1136 343 408 432 VSS nch l=0.04u w=0.4u
m1137 460 409 433 VSS nch l=0.04u w=0.4u
m1138 434 319 69365 VSS nch l=0.04u w=0.8u
m1139 FRAC[1] 410 435 VSS nch l=0.04u w=0.4u
m1140 343 411 436 VSS nch l=0.04u w=0.4u
m1141 463 4328 VSS VSS nch l=0.04u w=0.4u
m1142 464 4328 VSS VSS nch l=0.04u w=0.4u
m1143 465 4328 VSS VSS nch l=0.04u w=0.4u
m1144 466 4328 VSS VSS nch l=0.04u w=0.4u
m1145 69370 4328 426 VSS nch l=0.04u w=0.12u
m1146 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1147 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1148 VSS 479 69367 VSS nch l=0.04u w=0.12u
m1149 VSS 480 69368 VSS nch l=0.04u w=0.12u
m1150 455 336 69369 VSS nch l=0.04u w=0.8u
m1151 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1152 VSS 508 457 VSS nch l=0.04u w=0.4u
m1153 VSS 490 69370 VSS nch l=0.04u w=0.12u
m1154 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1155 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1156 VSS 467 467 VSS nch l=0.04u w=0.8u
m1157 VSS 470 470 VSS nch l=0.04u w=0.8u
m1158 479 413 VSS VSS nch l=0.04u w=0.4u
m1159 480 414 VSS VSS nch l=0.04u w=0.4u
m1160 69393 336 455 VSS nch l=0.04u w=0.8u
m1161 481 451 471 VSS nch l=0.04u w=0.4u
m1162 482 452 302 VSS nch l=0.04u w=0.4u
m1163 483 453 472 VSS nch l=0.04u w=0.4u
m1164 484 454 146 VSS nch l=0.04u w=0.4u
m1165 69394 521 456 VSS nch l=0.04u w=0.8u
m1166 69395 393 473 VSS nch l=0.04u w=0.8u
m1167 69396 394 475 VSS nch l=0.04u w=0.8u
m1168 490 426 VSS VSS nch l=0.04u w=0.4u
m1169 486 463 477 VSS nch l=0.04u w=0.4u
m1170 487 464 478 VSS nch l=0.04u w=0.4u
m1171 488 465 401 VSS nch l=0.04u w=0.4u
m1172 489 466 402 VSS nch l=0.04u w=0.4u
m1173 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1174 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1175 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1176 VSS 387 69393 VSS nch l=0.04u w=0.8u
m1177 69397 4328 481 VSS nch l=0.04u w=0.12u
m1178 69398 4328 482 VSS nch l=0.04u w=0.12u
m1179 69399 4328 483 VSS nch l=0.04u w=0.12u
m1180 69400 4328 484 VSS nch l=0.04u w=0.12u
m1181 VSS 2648 69394 VSS nch l=0.04u w=0.8u
m1182 VSS 508 485 VSS nch l=0.04u w=0.4u
m1183 VSS 206 69395 VSS nch l=0.04u w=0.8u
m1184 VSS 209 69396 VSS nch l=0.04u w=0.8u
m1185 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1186 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1187 69401 4328 486 VSS nch l=0.04u w=0.12u
m1188 69402 4328 487 VSS nch l=0.04u w=0.12u
m1189 69403 417 491 VSS nch l=0.04u w=0.8u
m1190 311 509 474 VSS nch l=0.04u w=0.4u
m1191 69404 419 492 VSS nch l=0.04u w=0.8u
m1192 69405 420 493 VSS nch l=0.04u w=0.8u
m1193 312 510 139 VSS nch l=0.04u w=0.4u
m1194 69406 422 494 VSS nch l=0.04u w=0.8u
m1195 69407 4328 488 VSS nch l=0.04u w=0.12u
m1196 69408 4328 489 VSS nch l=0.04u w=0.12u
m1197 69409 423 495 VSS nch l=0.04u w=0.8u
m1198 314 511 FRAC[23] VSS nch l=0.04u w=0.4u
m1199 69410 425 496 VSS nch l=0.04u w=0.8u
m1200 316 512 203 VSS nch l=0.04u w=0.4u
m1201 69411 428 497 VSS nch l=0.04u w=0.8u
m1202 69412 429 498 VSS nch l=0.04u w=0.8u
m1203 317 513 65 VSS nch l=0.04u w=0.4u
m1204 69413 431 499 VSS nch l=0.04u w=0.8u
m1205 69414 432 500 VSS nch l=0.04u w=0.8u
m1206 69415 433 501 VSS nch l=0.04u w=0.8u
m1207 319 514 FRAC[23] VSS nch l=0.04u w=0.4u
m1208 69416 435 502 VSS nch l=0.04u w=0.8u
m1209 69417 436 503 VSS nch l=0.04u w=0.8u
m1210 504 155 VSS VSS nch l=0.04u w=0.4u
m1211 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1212 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1213 505 4328 479 VSS nch l=0.04u w=0.4u
m1214 506 4328 480 VSS nch l=0.04u w=0.4u
m1215 VSS 516 69397 VSS nch l=0.04u w=0.12u
m1216 VSS 517 69398 VSS nch l=0.04u w=0.12u
m1217 VSS 518 69399 VSS nch l=0.04u w=0.12u
m1218 VSS 519 69400 VSS nch l=0.04u w=0.12u
m1219 69418 456 VSS VSS nch l=0.04u w=0.24u
m1220 VSS 523 69401 VSS nch l=0.04u w=0.12u
m1221 VSS 524 69402 VSS nch l=0.04u w=0.12u
m1222 VSS 218 69403 VSS nch l=0.04u w=0.8u
m1223 509 474 311 VSS nch l=0.04u w=0.4u
m1224 VSS 219 69404 VSS nch l=0.04u w=0.8u
m1225 VSS 220 69405 VSS nch l=0.04u w=0.8u
m1226 510 139 312 VSS nch l=0.04u w=0.4u
m1227 VSS 221 69406 VSS nch l=0.04u w=0.8u
m1228 VSS 526 69407 VSS nch l=0.04u w=0.12u
m1229 VSS 527 69408 VSS nch l=0.04u w=0.12u
m1230 VSS 222 69409 VSS nch l=0.04u w=0.8u
m1231 511 FRAC[23] 314 VSS nch l=0.04u w=0.4u
m1232 VSS 223 69410 VSS nch l=0.04u w=0.8u
m1233 507 4328 490 VSS nch l=0.04u w=0.4u
m1234 512 203 316 VSS nch l=0.04u w=0.4u
m1235 VSS 224 69411 VSS nch l=0.04u w=0.8u
m1236 VSS 225 69412 VSS nch l=0.04u w=0.8u
m1237 513 65 317 VSS nch l=0.04u w=0.4u
m1238 VSS 226 69413 VSS nch l=0.04u w=0.8u
m1239 VSS 227 69414 VSS nch l=0.04u w=0.8u
m1240 VSS 228 69415 VSS nch l=0.04u w=0.8u
m1241 514 FRAC[23] 319 VSS nch l=0.04u w=0.4u
m1242 VSS 229 69416 VSS nch l=0.04u w=0.8u
m1243 VSS 230 69417 VSS nch l=0.04u w=0.8u
m1244 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1245 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1246 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1247 69419 385 505 VSS nch l=0.04u w=0.12u
m1248 69420 386 506 VSS nch l=0.04u w=0.12u
m1249 516 481 VSS VSS nch l=0.04u w=0.4u
m1250 517 482 VSS VSS nch l=0.04u w=0.4u
m1251 518 483 VSS VSS nch l=0.04u w=0.4u
m1252 519 484 VSS VSS nch l=0.04u w=0.4u
m1253 520 76 VSS VSS nch l=0.04u w=0.4u
m1254 521 605 69418 VSS nch l=0.04u w=0.24u
m1255 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1256 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1257 69421 560 508 VSS nch l=0.04u w=0.8u
m1258 69422 473 VSS VSS nch l=0.04u w=0.8u
m1259 523 486 VSS VSS nch l=0.04u w=0.4u
m1260 524 487 VSS VSS nch l=0.04u w=0.4u
m1261 VSS 292 509 VSS nch l=0.04u w=0.4u
m1262 69423 475 VSS VSS nch l=0.04u w=0.8u
m1263 VSS 300 510 VSS nch l=0.04u w=0.4u
m1264 526 488 VSS VSS nch l=0.04u w=0.4u
m1265 527 489 VSS VSS nch l=0.04u w=0.4u
m1266 VSS 294 511 VSS nch l=0.04u w=0.4u
m1267 69424 390 507 VSS nch l=0.04u w=0.12u
m1268 VSS 347 512 VSS nch l=0.04u w=0.4u
m1269 VSS 203 513 VSS nch l=0.04u w=0.4u
m1270 VSS 205 514 VSS nch l=0.04u w=0.4u
m1271 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1272 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1273 69425 155 VSS VSS nch l=0.04u w=0.8u
m1274 VSS 548 69419 VSS nch l=0.04u w=0.12u
m1275 VSS 549 69420 VSS nch l=0.04u w=0.12u
m1276 VDDREF 561 521 VSS nch l=0.04u w=0.4u
m1277 VSS 764 69421 VSS nch l=0.04u w=0.8u
m1278 522 337 69422 VSS nch l=0.04u w=0.8u
m1279 525 338 69423 VSS nch l=0.04u w=0.8u
m1280 VSS 559 69424 VSS nch l=0.04u w=0.12u
m1281 69426 491 VSS VSS nch l=0.04u w=0.8u
m1282 69427 492 VSS VSS nch l=0.04u w=0.8u
m1283 69428 493 VSS VSS nch l=0.04u w=0.8u
m1284 69429 494 VSS VSS nch l=0.04u w=0.8u
m1285 69430 495 VSS VSS nch l=0.04u w=0.8u
m1286 69431 496 VSS VSS nch l=0.04u w=0.8u
m1287 69432 497 VSS VSS nch l=0.04u w=0.8u
m1288 69433 498 VSS VSS nch l=0.04u w=0.8u
m1289 69434 499 VSS VSS nch l=0.04u w=0.8u
m1290 69435 500 VSS VSS nch l=0.04u w=0.8u
m1291 69436 501 VSS VSS nch l=0.04u w=0.8u
m1292 69437 502 VSS VSS nch l=0.04u w=0.8u
m1293 69438 503 VSS VSS nch l=0.04u w=0.8u
m1294 528 FBDIV[1] 69425 VSS nch l=0.04u w=0.8u
m1295 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1296 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1297 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1298 548 505 VSS VSS nch l=0.04u w=0.4u
m1299 549 506 VSS VSS nch l=0.04u w=0.4u
m1300 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1301 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1302 550 4328 516 VSS nch l=0.04u w=0.4u
m1303 551 4328 517 VSS nch l=0.04u w=0.4u
m1304 552 4328 518 VSS nch l=0.04u w=0.4u
m1305 553 4328 519 VSS nch l=0.04u w=0.4u
m1306 554 520 455 VSS nch l=0.04u w=0.4u
m1307 559 507 VSS VSS nch l=0.04u w=0.4u
m1308 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1309 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1310 555 4328 523 VSS nch l=0.04u w=0.4u
m1311 556 4328 524 VSS nch l=0.04u w=0.4u
m1312 529 352 69426 VSS nch l=0.04u w=0.8u
m1313 69439 292 530 VSS nch l=0.04u w=0.8u
m1314 531 354 69427 VSS nch l=0.04u w=0.8u
m1315 532 355 69428 VSS nch l=0.04u w=0.8u
m1316 69440 300 533 VSS nch l=0.04u w=0.8u
m1317 534 357 69429 VSS nch l=0.04u w=0.8u
m1318 557 4328 526 VSS nch l=0.04u w=0.4u
m1319 558 4328 527 VSS nch l=0.04u w=0.4u
m1320 535 360 69430 VSS nch l=0.04u w=0.8u
m1321 69441 294 536 VSS nch l=0.04u w=0.8u
m1322 537 362 69431 VSS nch l=0.04u w=0.8u
m1323 69442 347 538 VSS nch l=0.04u w=0.8u
m1324 539 364 69432 VSS nch l=0.04u w=0.8u
m1325 540 365 69433 VSS nch l=0.04u w=0.8u
m1326 69443 203 541 VSS nch l=0.04u w=0.8u
m1327 542 367 69434 VSS nch l=0.04u w=0.8u
m1328 543 368 69435 VSS nch l=0.04u w=0.8u
m1329 544 369 69436 VSS nch l=0.04u w=0.8u
m1330 69444 205 545 VSS nch l=0.04u w=0.8u
m1331 546 371 69437 VSS nch l=0.04u w=0.8u
m1332 547 372 69438 VSS nch l=0.04u w=0.8u
m1333 69445 451 550 VSS nch l=0.04u w=0.12u
m1334 69446 452 551 VSS nch l=0.04u w=0.12u
m1335 69447 453 552 VSS nch l=0.04u w=0.12u
m1336 69448 454 553 VSS nch l=0.04u w=0.12u
m1337 69449 76 554 VSS nch l=0.04u w=0.12u
m1338 561 605 VSS VSS nch l=0.04u w=0.4u
m1339 VSS 594 560 VSS nch l=0.04u w=0.4u
m1340 562 393 VSS VSS nch l=0.04u w=0.4u
m1341 69450 463 555 VSS nch l=0.04u w=0.12u
m1342 69451 464 556 VSS nch l=0.04u w=0.12u
m1343 VSS 474 69439 VSS nch l=0.04u w=0.8u
m1344 563 394 VSS VSS nch l=0.04u w=0.4u
m1345 VSS 139 69440 VSS nch l=0.04u w=0.8u
m1346 69452 465 557 VSS nch l=0.04u w=0.12u
m1347 69453 466 558 VSS nch l=0.04u w=0.12u
m1348 VSS FRAC[23] 69441 VSS nch l=0.04u w=0.8u
m1349 VSS 203 69442 VSS nch l=0.04u w=0.8u
m1350 VSS 65 69443 VSS nch l=0.04u w=0.8u
m1351 VSS FRAC[23] 69444 VSS nch l=0.04u w=0.8u
m1352 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1353 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1354 69455 504 VSS VSS nch l=0.04u w=0.8u
m1355 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1356 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1357 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1358 565 4328 VSS VSS nch l=0.04u w=0.4u
m1359 566 4328 VSS VSS nch l=0.04u w=0.4u
m1360 VSS 589 69445 VSS nch l=0.04u w=0.12u
m1361 VSS 133 69446 VSS nch l=0.04u w=0.12u
m1362 VSS 590 69447 VSS nch l=0.04u w=0.12u
m1363 VSS 136 69448 VSS nch l=0.04u w=0.12u
m1364 VSS 591 69449 VSS nch l=0.04u w=0.12u
m1365 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1366 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1367 69456 485 VSS VSS nch l=0.04u w=0.12u
m1368 568 206 562 VSS nch l=0.04u w=0.4u
m1369 VSS 592 69450 VSS nch l=0.04u w=0.12u
m1370 VSS 438 69451 VSS nch l=0.04u w=0.12u
m1371 569 209 563 VSS nch l=0.04u w=0.4u
m1372 VSS 593 69452 VSS nch l=0.04u w=0.12u
m1373 VSS 442 69453 VSS nch l=0.04u w=0.12u
m1374 570 417 VSS VSS nch l=0.04u w=0.4u
m1375 572 419 VSS VSS nch l=0.04u w=0.4u
m1376 573 420 VSS VSS nch l=0.04u w=0.4u
m1377 575 422 VSS VSS nch l=0.04u w=0.4u
m1378 576 423 VSS VSS nch l=0.04u w=0.4u
m1379 578 425 VSS VSS nch l=0.04u w=0.4u
m1380 580 428 VSS VSS nch l=0.04u w=0.4u
m1381 581 429 VSS VSS nch l=0.04u w=0.4u
m1382 583 431 VSS VSS nch l=0.04u w=0.4u
m1383 584 432 VSS VSS nch l=0.04u w=0.4u
m1384 585 433 VSS VSS nch l=0.04u w=0.4u
m1385 587 435 VSS VSS nch l=0.04u w=0.4u
m1386 588 436 VSS VSS nch l=0.04u w=0.4u
m1387 564 559 69455 VSS nch l=0.04u w=0.8u
m1388 589 550 VSS VSS nch l=0.04u w=0.4u
m1389 133 551 VSS VSS nch l=0.04u w=0.4u
m1390 590 552 VSS VSS nch l=0.04u w=0.4u
m1391 136 553 VSS VSS nch l=0.04u w=0.4u
m1392 591 554 VSS VSS nch l=0.04u w=0.4u
m1393 VSS 605 567 VSS nch l=0.04u w=0.4u
m1394 594 753 69456 VSS nch l=0.04u w=0.12u
m1395 206 562 568 VSS nch l=0.04u w=0.4u
m1396 592 555 VSS VSS nch l=0.04u w=0.4u
m1397 438 556 VSS VSS nch l=0.04u w=0.4u
m1398 VSS 340 VSS VSS nch l=0.26u w=0.8u
m1399 209 563 569 VSS nch l=0.04u w=0.4u
m1400 593 557 VSS VSS nch l=0.04u w=0.4u
m1401 442 558 VSS VSS nch l=0.04u w=0.4u
m1402 VSS 342 VSS VSS nch l=0.26u w=0.8u
m1403 595 218 570 VSS nch l=0.04u w=0.4u
m1404 478 219 572 VSS nch l=0.04u w=0.4u
m1405 596 220 573 VSS nch l=0.04u w=0.4u
m1406 598 221 575 VSS nch l=0.04u w=0.4u
m1407 439 222 576 VSS nch l=0.04u w=0.4u
m1408 440 223 578 VSS nch l=0.04u w=0.4u
m1409 412 224 580 VSS nch l=0.04u w=0.4u
m1410 601 225 581 VSS nch l=0.04u w=0.4u
m1411 262 226 583 VSS nch l=0.04u w=0.4u
m1412 462 227 584 VSS nch l=0.04u w=0.4u
m1413 444 228 585 VSS nch l=0.04u w=0.4u
m1414 264 229 587 VSS nch l=0.04u w=0.4u
m1415 460 230 588 VSS nch l=0.04u w=0.4u
m1416 VSS 345 VSS VSS nch l=0.26u w=0.8u
m1417 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1418 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1419 602 565 548 VSS nch l=0.04u w=0.4u
m1420 603 566 549 VSS nch l=0.04u w=0.4u
m1421 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1422 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1423 604 76 594 VSS nch l=0.04u w=0.4u
m1424 606 607 VSS VSS nch l=0.04u w=0.8u
m1425 608 609 VSS VSS nch l=0.04u w=0.8u
m1426 218 570 595 VSS nch l=0.04u w=0.4u
m1427 219 572 478 VSS nch l=0.04u w=0.4u
m1428 220 573 596 VSS nch l=0.04u w=0.4u
m1429 221 575 598 VSS nch l=0.04u w=0.4u
m1430 222 576 439 VSS nch l=0.04u w=0.4u
m1431 223 578 440 VSS nch l=0.04u w=0.4u
m1432 224 580 412 VSS nch l=0.04u w=0.4u
m1433 225 581 601 VSS nch l=0.04u w=0.4u
m1434 226 583 262 VSS nch l=0.04u w=0.4u
m1435 227 584 462 VSS nch l=0.04u w=0.4u
m1436 228 585 444 VSS nch l=0.04u w=0.4u
m1437 229 587 264 VSS nch l=0.04u w=0.4u
m1438 230 588 460 VSS nch l=0.04u w=0.4u
m1439 477 624 571 VSS nch l=0.04u w=0.4u
m1440 597 625 574 VSS nch l=0.04u w=0.4u
m1441 599 626 577 VSS nch l=0.04u w=0.4u
m1442 600 627 579 VSS nch l=0.04u w=0.4u
m1443 62 628 582 VSS nch l=0.04u w=0.4u
m1444 64 629 586 VSS nch l=0.04u w=0.4u
m1445 69466 564 VSS VSS nch l=0.04u w=0.8u
m1446 617 618 VSS VSS nch l=0.04u w=0.8u
m1447 69473 4328 602 VSS nch l=0.04u w=0.12u
m1448 69474 4328 603 VSS nch l=0.04u w=0.12u
m1449 620 4328 VSS VSS nch l=0.04u w=0.4u
m1450 621 4328 VSS VSS nch l=0.04u w=0.4u
m1451 622 4328 VSS VSS nch l=0.04u w=0.4u
m1452 623 4328 VSS VSS nch l=0.04u w=0.4u
m1453 619 76 591 VSS nch l=0.04u w=0.4u
m1454 69475 652 605 VSS nch l=0.04u w=0.8u
m1455 624 571 477 VSS nch l=0.04u w=0.4u
m1456 625 574 597 VSS nch l=0.04u w=0.4u
m1457 626 577 599 VSS nch l=0.04u w=0.4u
m1458 627 579 600 VSS nch l=0.04u w=0.4u
m1459 628 582 62 VSS nch l=0.04u w=0.4u
m1460 629 586 64 VSS nch l=0.04u w=0.4u
m1461 616 528 69466 VSS nch l=0.04u w=0.8u
m1462 VSS 380 VSS VSS nch l=0.26u w=0.8u
m1463 VSS 383 VSS VSS nch l=0.26u w=0.8u
m1464 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1465 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1466 VSS 646 69473 VSS nch l=0.04u w=0.12u
m1467 VSS 647 69474 VSS nch l=0.04u w=0.12u
m1468 69494 520 619 VSS nch l=0.04u w=0.12u
m1469 VSS 2648 69475 VSS nch l=0.04u w=0.8u
m1470 69495 675 604 VSS nch l=0.04u w=0.8u
m1471 69498 710 VSS VSS nch l=0.04u w=0.8u
m1472 VSS 610 624 VSS nch l=0.04u w=0.4u
m1473 69499 672 VSS VSS nch l=0.04u w=0.8u
m1474 VSS 611 625 VSS nch l=0.04u w=0.4u
m1475 VSS 612 626 VSS nch l=0.04u w=0.4u
m1476 VSS 613 627 VSS nch l=0.04u w=0.4u
m1477 VSS 614 628 VSS nch l=0.04u w=0.4u
m1478 VSS 615 629 VSS nch l=0.04u w=0.4u
m1479 VSS 630 630 VSS nch l=0.04u w=0.8u
m1480 643 642 VSS VSS nch l=0.04u w=0.8u
m1481 644 645 VSS VSS nch l=0.04u w=0.8u
m1482 646 602 VSS VSS nch l=0.04u w=0.4u
m1483 647 603 VSS VSS nch l=0.04u w=0.4u
m1484 VSS 259 69494 VSS nch l=0.04u w=0.12u
m1485 648 620 633 VSS nch l=0.04u w=0.4u
m1486 649 621 601 VSS nch l=0.04u w=0.4u
m1487 650 622 634 VSS nch l=0.04u w=0.4u
m1488 651 623 444 VSS nch l=0.04u w=0.4u
m1489 VSS 764 69495 VSS nch l=0.04u w=0.8u
m1490 635 688 69498 VSS nch l=0.04u w=0.8u
m1491 636 593 69499 VSS nch l=0.04u w=0.8u
m1492 VSS 637 637 VSS nch l=0.04u w=0.8u
m1493 69501 754 VSS VSS nch l=0.04u w=0.8u
m1494 69502 736 VSS VSS nch l=0.04u w=0.8u
m1495 69503 139 VSS VSS nch l=0.04u w=0.8u
m1496 69504 755 VSS VSS nch l=0.04u w=0.8u
m1497 69505 2616 VSS VSS nch l=0.04u w=0.8u
m1498 69506 2616 VSS VSS nch l=0.04u w=0.8u
m1499 VSS 639 639 VSS nch l=0.04u w=0.8u
m1500 69507 756 VSS VSS nch l=0.04u w=0.8u
m1501 69508 FRAC[2] VSS VSS nch l=0.04u w=0.8u
m1502 VSS 704 641 VSS nch l=0.04u w=0.4u
m1503 69509 737 VSS VSS nch l=0.04u w=0.8u
m1504 69510 758 VSS VSS nch l=0.04u w=0.8u
m1505 69511 634 VSS VSS nch l=0.04u w=0.8u
m1506 69512 641 VSS VSS nch l=0.04u w=0.8u
m1507 69513 756 VSS VSS nch l=0.04u w=0.8u
m1508 69514 FRAC[2] VSS VSS nch l=0.04u w=0.8u
m1509 69515 641 VSS VSS nch l=0.04u w=0.8u
m1510 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1511 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1512 259 619 VSS VSS nch l=0.04u w=0.4u
m1513 69516 4328 648 VSS nch l=0.04u w=0.12u
m1514 69517 4328 649 VSS nch l=0.04u w=0.12u
m1515 69518 4328 650 VSS nch l=0.04u w=0.12u
m1516 69519 4328 651 VSS nch l=0.04u w=0.12u
m1517 69520 604 VSS VSS nch l=0.04u w=0.24u
m1518 VSS 685 652 VSS nch l=0.04u w=0.4u
m1519 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1520 653 731 69501 VSS nch l=0.04u w=0.8u
m1521 69522 823 274 VSS nch l=0.04u w=0.8u
m1522 654 732 69502 VSS nch l=0.04u w=0.8u
m1523 655 733 69503 VSS nch l=0.04u w=0.8u
m1524 69523 826 277 VSS nch l=0.04u w=0.8u
m1525 656 734 69504 VSS nch l=0.04u w=0.8u
m1526 657 893 69505 VSS nch l=0.04u w=0.8u
m1527 658 894 69506 VSS nch l=0.04u w=0.8u
m1528 659 735 69507 VSS nch l=0.04u w=0.8u
m1529 69524 829 280 VSS nch l=0.04u w=0.8u
m1530 660 736 69508 VSS nch l=0.04u w=0.8u
m1531 69525 831 282 VSS nch l=0.04u w=0.8u
m1532 661 131 69509 VSS nch l=0.04u w=0.8u
m1533 662 737 69510 VSS nch l=0.04u w=0.8u
m1534 69526 834 285 VSS nch l=0.04u w=0.8u
m1535 663 738 69511 VSS nch l=0.04u w=0.8u
m1536 664 739 69512 VSS nch l=0.04u w=0.8u
m1537 665 740 69513 VSS nch l=0.04u w=0.8u
m1538 69527 838 289 VSS nch l=0.04u w=0.8u
m1539 666 741 69514 VSS nch l=0.04u w=0.8u
m1540 667 FBDIV[2] 69515 VSS nch l=0.04u w=0.8u
m1541 VSS 669 669 VSS nch l=0.04u w=0.8u
m1542 VSS 670 670 VSS nch l=0.04u w=0.8u
m1543 673 4328 646 VSS nch l=0.04u w=0.4u
m1544 674 4328 647 VSS nch l=0.04u w=0.4u
m1545 VSS 679 69516 VSS nch l=0.04u w=0.12u
m1546 VSS 680 69517 VSS nch l=0.04u w=0.12u
m1547 VSS 681 69518 VSS nch l=0.04u w=0.12u
m1548 VSS 682 69519 VSS nch l=0.04u w=0.12u
m1549 675 76 69520 VSS nch l=0.04u w=0.24u
m1550 69529 567 VSS VSS nch l=0.04u w=0.12u
m1551 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1552 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1553 676 688 VSS VSS nch l=0.04u w=0.4u
m1554 VSS 712 69522 VSS nch l=0.04u w=0.8u
m1555 677 593 VSS VSS nch l=0.04u w=0.4u
m1556 VSS 715 69523 VSS nch l=0.04u w=0.8u
m1557 VSS 718 69524 VSS nch l=0.04u w=0.8u
m1558 VSS 721 69525 VSS nch l=0.04u w=0.8u
m1559 VSS 724 69526 VSS nch l=0.04u w=0.8u
m1560 VSS 728 69527 VSS nch l=0.04u w=0.8u
m1561 678 4328 VSS VSS nch l=0.04u w=0.4u
m1562 VSS 2197 672 VSS nch l=0.04u w=0.4u
m1563 VSS 468 VSS VSS nch l=0.26u w=0.8u
m1564 VSS 469 VSS VSS nch l=0.26u w=0.8u
m1565 69532 565 673 VSS nch l=0.04u w=0.12u
m1566 69533 566 674 VSS nch l=0.04u w=0.12u
m1567 679 648 VSS VSS nch l=0.04u w=0.4u
m1568 680 649 VSS VSS nch l=0.04u w=0.4u
m1569 681 650 VSS VSS nch l=0.04u w=0.4u
m1570 682 651 VSS VSS nch l=0.04u w=0.4u
m1571 683 259 VSS VSS nch l=0.04u w=0.4u
m1572 684 753 675 VSS nch l=0.04u w=0.4u
m1573 685 847 69529 VSS nch l=0.04u w=0.12u
m1574 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1575 686 710 676 VSS nch l=0.04u w=0.4u
m1576 687 672 677 VSS nch l=0.04u w=0.4u
m1577 689 731 VSS VSS nch l=0.04u w=0.4u
m1578 690 732 VSS VSS nch l=0.04u w=0.4u
m1579 691 733 VSS VSS nch l=0.04u w=0.4u
m1580 692 734 VSS VSS nch l=0.04u w=0.4u
m1581 693 657 VSS VSS nch l=0.04u w=0.4u
m1582 694 658 VSS VSS nch l=0.04u w=0.4u
m1583 695 735 VSS VSS nch l=0.04u w=0.4u
m1584 696 736 VSS VSS nch l=0.04u w=0.4u
m1585 697 131 VSS VSS nch l=0.04u w=0.4u
m1586 698 737 VSS VSS nch l=0.04u w=0.4u
m1587 699 738 VSS VSS nch l=0.04u w=0.4u
m1588 700 739 VSS VSS nch l=0.04u w=0.4u
m1589 701 740 VSS VSS nch l=0.04u w=0.4u
m1590 702 741 VSS VSS nch l=0.04u w=0.4u
m1591 703 FBDIV[2] VSS VSS nch l=0.04u w=0.4u
m1592 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1593 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1594 705 706 VSS VSS nch l=0.04u w=0.8u
m1595 708 707 VSS VSS nch l=0.04u w=0.8u
m1596 VSS 747 69532 VSS nch l=0.04u w=0.12u
m1597 VSS 748 69533 VSS nch l=0.04u w=0.12u
m1598 VSS 259 683 VSS nch l=0.04u w=0.4u
m1599 709 886 685 VSS nch l=0.04u w=0.4u
m1600 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1601 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1602 710 676 686 VSS nch l=0.04u w=0.4u
m1603 672 677 687 VSS nch l=0.04u w=0.4u
m1604 711 754 689 VSS nch l=0.04u w=0.4u
m1605 69534 571 VSS VSS nch l=0.04u w=0.8u
m1606 713 736 690 VSS nch l=0.04u w=0.4u
m1607 714 139 691 VSS nch l=0.04u w=0.4u
m1608 69535 574 VSS VSS nch l=0.04u w=0.8u
m1609 716 755 692 VSS nch l=0.04u w=0.4u
m1610 717 756 695 VSS nch l=0.04u w=0.4u
m1611 69536 577 VSS VSS nch l=0.04u w=0.8u
m1612 719 FRAC[2] 696 VSS nch l=0.04u w=0.4u
m1613 69537 579 VSS VSS nch l=0.04u w=0.8u
m1614 722 737 697 VSS nch l=0.04u w=0.4u
m1615 723 758 698 VSS nch l=0.04u w=0.4u
m1616 69538 582 VSS VSS nch l=0.04u w=0.8u
m1617 725 634 699 VSS nch l=0.04u w=0.4u
m1618 726 641 700 VSS nch l=0.04u w=0.4u
m1619 727 756 701 VSS nch l=0.04u w=0.4u
m1620 69539 586 VSS VSS nch l=0.04u w=0.8u
m1621 729 FRAC[2] 702 VSS nch l=0.04u w=0.4u
m1622 730 641 703 VSS nch l=0.04u w=0.4u
m1623 720 678 704 VSS nch l=0.04u w=0.4u
m1624 747 673 VSS VSS nch l=0.04u w=0.4u
m1625 748 674 VSS VSS nch l=0.04u w=0.4u
m1626 749 4328 679 VSS nch l=0.04u w=0.4u
m1627 750 4328 680 VSS nch l=0.04u w=0.4u
m1628 751 4328 681 VSS nch l=0.04u w=0.4u
m1629 752 4328 682 VSS nch l=0.04u w=0.4u
m1630 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1631 753 76 VSS VSS nch l=0.04u w=0.4u
m1632 754 689 711 VSS nch l=0.04u w=0.4u
m1633 712 610 69534 VSS nch l=0.04u w=0.8u
m1634 736 690 713 VSS nch l=0.04u w=0.4u
m1635 139 691 714 VSS nch l=0.04u w=0.4u
m1636 715 611 69535 VSS nch l=0.04u w=0.8u
m1637 755 692 716 VSS nch l=0.04u w=0.4u
m1638 756 695 717 VSS nch l=0.04u w=0.4u
m1639 718 612 69536 VSS nch l=0.04u w=0.8u
m1640 FRAC[2] 696 719 VSS nch l=0.04u w=0.4u
m1641 721 613 69537 VSS nch l=0.04u w=0.8u
m1642 737 697 722 VSS nch l=0.04u w=0.4u
m1643 758 698 723 VSS nch l=0.04u w=0.4u
m1644 724 614 69538 VSS nch l=0.04u w=0.8u
m1645 634 699 725 VSS nch l=0.04u w=0.4u
m1646 641 700 726 VSS nch l=0.04u w=0.4u
m1647 756 701 727 VSS nch l=0.04u w=0.4u
m1648 728 615 69539 VSS nch l=0.04u w=0.8u
m1649 FRAC[2] 702 729 VSS nch l=0.04u w=0.4u
m1650 641 703 730 VSS nch l=0.04u w=0.4u
m1651 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1652 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1653 759 4328 VSS VSS nch l=0.04u w=0.4u
m1654 760 4328 VSS VSS nch l=0.04u w=0.4u
m1655 761 4328 VSS VSS nch l=0.04u w=0.4u
m1656 762 4328 VSS VSS nch l=0.04u w=0.4u
m1657 69541 4328 720 VSS nch l=0.04u w=0.12u
m1658 VSS 743 743 VSS nch l=0.04u w=0.8u
m1659 VSS 746 746 VSS nch l=0.04u w=0.8u
m1660 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1661 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1662 69545 620 749 VSS nch l=0.04u w=0.12u
m1663 69546 621 750 VSS nch l=0.04u w=0.12u
m1664 69547 622 751 VSS nch l=0.04u w=0.12u
m1665 69548 623 752 VSS nch l=0.04u w=0.12u
m1666 763 683 VSS VSS nch l=0.04u w=0.4u
m1667 69549 798 709 VSS nch l=0.04u w=0.8u
m1668 VSS 778 69541 VSS nch l=0.04u w=0.12u
m1669 771 4328 VSS VSS nch l=0.04u w=0.4u
m1670 772 4328 VSS VSS nch l=0.04u w=0.4u
m1671 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1672 VSS 738 69545 VSS nch l=0.04u w=0.12u
m1673 VSS 443 69546 VSS nch l=0.04u w=0.12u
m1674 VSS 741 69547 VSS nch l=0.04u w=0.12u
m1675 VSS 445 69548 VSS nch l=0.04u w=0.12u
m1676 VSS 2648 69549 VSS nch l=0.04u w=0.8u
m1677 VSS 236 764 VSS nch l=0.04u w=0.4u
m1678 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1679 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1680 69569 686 765 VSS nch l=0.04u w=0.8u
m1681 69570 687 767 VSS nch l=0.04u w=0.8u
m1682 778 720 VSS VSS nch l=0.04u w=0.4u
m1683 774 759 769 VSS nch l=0.04u w=0.4u
m1684 775 760 770 VSS nch l=0.04u w=0.4u
m1685 776 761 693 VSS nch l=0.04u w=0.4u
m1686 777 762 694 VSS nch l=0.04u w=0.4u
m1687 VSS 744 VSS VSS nch l=0.26u w=0.8u
m1688 VSS 745 VSS VSS nch l=0.26u w=0.8u
m1689 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1690 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1691 738 749 VSS VSS nch l=0.04u w=0.4u
m1692 443 750 VSS VSS nch l=0.04u w=0.4u
m1693 741 751 VSS VSS nch l=0.04u w=0.4u
m1694 445 752 VSS VSS nch l=0.04u w=0.4u
m1695 792 763 VSS VSS nch l=0.04u w=0.4u
m1696 69571 709 VSS VSS nch l=0.04u w=0.24u
m1697 VSS 522 69569 VSS nch l=0.04u w=0.8u
m1698 VSS 525 69570 VSS nch l=0.04u w=0.8u
m1699 69572 4328 774 VSS nch l=0.04u w=0.12u
m1700 69573 4328 775 VSS nch l=0.04u w=0.12u
m1701 69574 711 779 VSS nch l=0.04u w=0.8u
m1702 610 800 766 VSS nch l=0.04u w=0.4u
m1703 69575 713 780 VSS nch l=0.04u w=0.8u
m1704 69576 714 781 VSS nch l=0.04u w=0.8u
m1705 611 801 139 VSS nch l=0.04u w=0.4u
m1706 69577 716 782 VSS nch l=0.04u w=0.8u
m1707 69578 4328 776 VSS nch l=0.04u w=0.12u
m1708 69579 4328 777 VSS nch l=0.04u w=0.12u
m1709 69580 717 783 VSS nch l=0.04u w=0.8u
m1710 612 802 FRAC[22] VSS nch l=0.04u w=0.4u
m1711 69581 719 784 VSS nch l=0.04u w=0.8u
m1712 613 803 202 VSS nch l=0.04u w=0.4u
m1713 69582 722 785 VSS nch l=0.04u w=0.8u
m1714 69583 723 786 VSS nch l=0.04u w=0.8u
m1715 614 804 64 VSS nch l=0.04u w=0.4u
m1716 69584 725 787 VSS nch l=0.04u w=0.8u
m1717 69585 726 788 VSS nch l=0.04u w=0.8u
m1718 69586 727 789 VSS nch l=0.04u w=0.8u
m1719 615 805 FRAC[22] VSS nch l=0.04u w=0.4u
m1720 69587 729 790 VSS nch l=0.04u w=0.8u
m1721 69588 730 791 VSS nch l=0.04u w=0.8u
m1722 794 155 VSS VSS nch l=0.04u w=0.4u
m1723 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1724 795 771 747 VSS nch l=0.04u w=0.4u
m1725 796 772 748 VSS nch l=0.04u w=0.4u
m1726 798 886 69571 VSS nch l=0.04u w=0.24u
m1727 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1728 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1729 69589 683 684 VSS nch l=0.04u w=0.8u
m1730 VSS 744 VSS VSS nch l=0.26u w=0.8u
m1731 VSS 745 VSS VSS nch l=0.26u w=0.8u
m1732 VSS 812 69572 VSS nch l=0.04u w=0.12u
m1733 VSS 813 69573 VSS nch l=0.04u w=0.12u
m1734 VSS 529 69574 VSS nch l=0.04u w=0.8u
m1735 800 766 610 VSS nch l=0.04u w=0.4u
m1736 VSS 531 69575 VSS nch l=0.04u w=0.8u
m1737 VSS 532 69576 VSS nch l=0.04u w=0.8u
m1738 801 139 611 VSS nch l=0.04u w=0.4u
m1739 VSS 534 69577 VSS nch l=0.04u w=0.8u
m1740 VSS 815 69578 VSS nch l=0.04u w=0.12u
m1741 VSS 816 69579 VSS nch l=0.04u w=0.12u
m1742 VSS 535 69580 VSS nch l=0.04u w=0.8u
m1743 802 FRAC[22] 612 VSS nch l=0.04u w=0.4u
m1744 VSS 537 69581 VSS nch l=0.04u w=0.8u
m1745 799 4328 778 VSS nch l=0.04u w=0.4u
m1746 803 202 613 VSS nch l=0.04u w=0.4u
m1747 VSS 539 69582 VSS nch l=0.04u w=0.8u
m1748 VSS 540 69583 VSS nch l=0.04u w=0.8u
m1749 804 64 614 VSS nch l=0.04u w=0.4u
m1750 VSS 542 69584 VSS nch l=0.04u w=0.8u
m1751 VSS 543 69585 VSS nch l=0.04u w=0.8u
m1752 VSS 544 69586 VSS nch l=0.04u w=0.8u
m1753 805 FRAC[22] 615 VSS nch l=0.04u w=0.4u
m1754 VSS 546 69587 VSS nch l=0.04u w=0.8u
m1755 VSS 547 69588 VSS nch l=0.04u w=0.8u
m1756 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1757 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1758 69590 4328 795 VSS nch l=0.04u w=0.12u
m1759 69591 4328 796 VSS nch l=0.04u w=0.12u
m1760 806 4328 VSS VSS nch l=0.04u w=0.4u
m1761 807 4328 VSS VSS nch l=0.04u w=0.4u
m1762 808 4328 VSS VSS nch l=0.04u w=0.4u
m1763 809 4328 VSS VSS nch l=0.04u w=0.4u
m1764 605 847 798 VSS nch l=0.04u w=0.4u
m1765 797 810 763 VSS nch l=0.04u w=0.4u
m1766 VSS 821 69589 VSS nch l=0.04u w=0.8u
m1767 69592 765 VSS VSS nch l=0.04u w=0.8u
m1768 812 774 VSS VSS nch l=0.04u w=0.4u
m1769 813 775 VSS VSS nch l=0.04u w=0.4u
m1770 VSS 592 800 VSS nch l=0.04u w=0.4u
m1771 69593 767 VSS VSS nch l=0.04u w=0.8u
m1772 VSS 599 801 VSS nch l=0.04u w=0.4u
m1773 815 776 VSS VSS nch l=0.04u w=0.4u
m1774 816 777 VSS VSS nch l=0.04u w=0.4u
m1775 VSS 593 802 VSS nch l=0.04u w=0.4u
m1776 69594 678 799 VSS nch l=0.04u w=0.12u
m1777 VSS 793 803 VSS nch l=0.04u w=0.4u
m1778 VSS 202 804 VSS nch l=0.04u w=0.4u
m1779 VSS 204 805 VSS nch l=0.04u w=0.4u
m1780 69595 155 VSS VSS nch l=0.04u w=0.8u
m1781 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1782 VSS 841 69590 VSS nch l=0.04u w=0.12u
m1783 VSS 842 69591 VSS nch l=0.04u w=0.12u
m1784 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1785 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1786 810 763 797 VSS nch l=0.04u w=0.4u
m1787 VSS 744 VSS VSS nch l=0.26u w=0.8u
m1788 VSS 745 VSS VSS nch l=0.26u w=0.8u
m1789 811 635 69592 VSS nch l=0.04u w=0.8u
m1790 814 636 69593 VSS nch l=0.04u w=0.8u
m1791 VSS 852 69594 VSS nch l=0.04u w=0.12u
m1792 69596 779 VSS VSS nch l=0.04u w=0.8u
m1793 69597 780 VSS VSS nch l=0.04u w=0.8u
m1794 69598 781 VSS VSS nch l=0.04u w=0.8u
m1795 69599 782 VSS VSS nch l=0.04u w=0.8u
m1796 69600 783 VSS VSS nch l=0.04u w=0.8u
m1797 69601 784 VSS VSS nch l=0.04u w=0.8u
m1798 69602 785 VSS VSS nch l=0.04u w=0.8u
m1799 69603 786 VSS VSS nch l=0.04u w=0.8u
m1800 69604 787 VSS VSS nch l=0.04u w=0.8u
m1801 69605 788 VSS VSS nch l=0.04u w=0.8u
m1802 69606 789 VSS VSS nch l=0.04u w=0.8u
m1803 69607 790 VSS VSS nch l=0.04u w=0.8u
m1804 69608 791 VSS VSS nch l=0.04u w=0.8u
m1805 817 FBDIV[2] 69595 VSS nch l=0.04u w=0.8u
m1806 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1807 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1808 841 795 VSS VSS nch l=0.04u w=0.4u
m1809 842 796 VSS VSS nch l=0.04u w=0.4u
m1810 843 806 818 VSS nch l=0.04u w=0.4u
m1811 844 807 819 VSS nch l=0.04u w=0.4u
m1812 845 808 820 VSS nch l=0.04u w=0.4u
m1813 846 809 739 VSS nch l=0.04u w=0.4u
m1814 847 886 VSS VSS nch l=0.04u w=0.4u
m1815 VSS 855 821 VSS nch l=0.04u w=0.4u
m1816 852 799 VSS VSS nch l=0.04u w=0.4u
m1817 848 4328 812 VSS nch l=0.04u w=0.4u
m1818 849 4328 813 VSS nch l=0.04u w=0.4u
m1819 822 653 69596 VSS nch l=0.04u w=0.8u
m1820 69609 592 823 VSS nch l=0.04u w=0.8u
m1821 824 654 69597 VSS nch l=0.04u w=0.8u
m1822 825 655 69598 VSS nch l=0.04u w=0.8u
m1823 69610 599 826 VSS nch l=0.04u w=0.8u
m1824 827 656 69599 VSS nch l=0.04u w=0.8u
m1825 850 4328 815 VSS nch l=0.04u w=0.4u
m1826 851 4328 816 VSS nch l=0.04u w=0.4u
m1827 828 659 69600 VSS nch l=0.04u w=0.8u
m1828 69611 593 829 VSS nch l=0.04u w=0.8u
m1829 830 660 69601 VSS nch l=0.04u w=0.8u
m1830 69612 793 831 VSS nch l=0.04u w=0.8u
m1831 832 661 69602 VSS nch l=0.04u w=0.8u
m1832 833 662 69603 VSS nch l=0.04u w=0.8u
m1833 69613 202 834 VSS nch l=0.04u w=0.8u
m1834 835 663 69604 VSS nch l=0.04u w=0.8u
m1835 836 664 69605 VSS nch l=0.04u w=0.8u
m1836 837 665 69606 VSS nch l=0.04u w=0.8u
m1837 69614 204 838 VSS nch l=0.04u w=0.8u
m1838 839 666 69607 VSS nch l=0.04u w=0.8u
m1839 840 667 69608 VSS nch l=0.04u w=0.8u
m1840 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1841 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1842 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1843 69615 4328 843 VSS nch l=0.04u w=0.12u
m1844 69616 4328 844 VSS nch l=0.04u w=0.12u
m1845 69617 4328 845 VSS nch l=0.04u w=0.12u
m1846 69618 4328 846 VSS nch l=0.04u w=0.12u
m1847 VSS 744 VSS VSS nch l=0.26u w=0.8u
m1848 VSS 745 VSS VSS nch l=0.26u w=0.8u
m1849 853 377 VSS VSS nch l=0.04u w=0.4u
m1850 856 686 VSS VSS nch l=0.04u w=0.4u
m1851 69619 759 848 VSS nch l=0.04u w=0.12u
m1852 69620 760 849 VSS nch l=0.04u w=0.12u
m1853 VSS 766 69609 VSS nch l=0.04u w=0.8u
m1854 857 687 VSS VSS nch l=0.04u w=0.4u
m1855 VSS 139 69610 VSS nch l=0.04u w=0.8u
m1856 69621 761 850 VSS nch l=0.04u w=0.12u
m1857 69622 762 851 VSS nch l=0.04u w=0.12u
m1858 VSS FRAC[22] 69611 VSS nch l=0.04u w=0.8u
m1859 VSS 202 69612 VSS nch l=0.04u w=0.8u
m1860 VSS 64 69613 VSS nch l=0.04u w=0.8u
m1861 VSS FRAC[22] 69614 VSS nch l=0.04u w=0.8u
m1862 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1863 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1864 69624 794 VSS VSS nch l=0.04u w=0.8u
m1865 859 4328 841 VSS nch l=0.04u w=0.4u
m1866 860 4328 842 VSS nch l=0.04u w=0.4u
m1867 VSS 881 69615 VSS nch l=0.04u w=0.12u
m1868 VSS 882 69616 VSS nch l=0.04u w=0.12u
m1869 VSS 883 69617 VSS nch l=0.04u w=0.12u
m1870 VSS 884 69618 VSS nch l=0.04u w=0.12u
m1871 VSS 886 854 VSS nch l=0.04u w=0.4u
m1872 69625 1000 855 VSS nch l=0.04u w=0.8u
m1873 861 522 856 VSS nch l=0.04u w=0.4u
m1874 VSS 888 69619 VSS nch l=0.04u w=0.12u
m1875 VSS 732 69620 VSS nch l=0.04u w=0.12u
m1876 766 525 857 VSS nch l=0.04u w=0.4u
m1877 VSS 398 69621 VSS nch l=0.04u w=0.12u
m1878 VSS 736 69622 VSS nch l=0.04u w=0.12u
m1879 VSS 631 VSS VSS nch l=0.26u w=0.8u
m1880 862 711 VSS VSS nch l=0.04u w=0.4u
m1881 864 713 VSS VSS nch l=0.04u w=0.4u
m1882 865 714 VSS VSS nch l=0.04u w=0.4u
m1883 867 716 VSS VSS nch l=0.04u w=0.4u
m1884 868 717 VSS VSS nch l=0.04u w=0.4u
m1885 870 719 VSS VSS nch l=0.04u w=0.4u
m1886 872 722 VSS VSS nch l=0.04u w=0.4u
m1887 873 723 VSS VSS nch l=0.04u w=0.4u
m1888 875 725 VSS VSS nch l=0.04u w=0.4u
m1889 876 726 VSS VSS nch l=0.04u w=0.4u
m1890 877 727 VSS VSS nch l=0.04u w=0.4u
m1891 879 729 VSS VSS nch l=0.04u w=0.4u
m1892 880 730 VSS VSS nch l=0.04u w=0.4u
m1893 858 852 69624 VSS nch l=0.04u w=0.8u
m1894 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1895 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1896 69632 771 859 VSS nch l=0.04u w=0.12u
m1897 69633 772 860 VSS nch l=0.04u w=0.12u
m1898 881 843 VSS VSS nch l=0.04u w=0.4u
m1899 882 844 VSS VSS nch l=0.04u w=0.4u
m1900 883 845 VSS VSS nch l=0.04u w=0.4u
m1901 884 846 VSS VSS nch l=0.04u w=0.4u
m1902 VSS 744 VSS VSS nch l=0.26u w=0.8u
m1903 VSS 745 VSS VSS nch l=0.26u w=0.8u
m1904 69634 377 VSS VSS nch l=0.04u w=0.8u
m1905 69635 918 69625 VSS nch l=0.04u w=0.8u
m1906 522 856 861 VSS nch l=0.04u w=0.4u
m1907 888 848 VSS VSS nch l=0.04u w=0.4u
m1908 732 849 VSS VSS nch l=0.04u w=0.4u
m1909 VSS 638 VSS VSS nch l=0.26u w=0.8u
m1910 525 857 766 VSS nch l=0.04u w=0.4u
m1911 398 850 VSS VSS nch l=0.04u w=0.4u
m1912 736 851 VSS VSS nch l=0.04u w=0.4u
m1913 VSS 640 VSS VSS nch l=0.26u w=0.8u
m1914 889 890 VSS VSS nch l=0.04u w=0.8u
m1915 891 529 862 VSS nch l=0.04u w=0.4u
m1916 770 531 864 VSS nch l=0.04u w=0.4u
m1917 892 532 865 VSS nch l=0.04u w=0.4u
m1918 894 534 867 VSS nch l=0.04u w=0.4u
m1919 733 535 868 VSS nch l=0.04u w=0.4u
m1920 734 537 870 VSS nch l=0.04u w=0.4u
m1921 704 539 872 VSS nch l=0.04u w=0.4u
m1922 819 540 873 VSS nch l=0.04u w=0.4u
m1923 633 542 875 VSS nch l=0.04u w=0.4u
m1924 758 543 876 VSS nch l=0.04u w=0.4u
m1925 739 544 877 VSS nch l=0.04u w=0.4u
m1926 634 546 879 VSS nch l=0.04u w=0.4u
m1927 756 547 880 VSS nch l=0.04u w=0.4u
m1928 VSS 912 69632 VSS nch l=0.04u w=0.12u
m1929 VSS 913 69633 VSS nch l=0.04u w=0.12u
m1930 898 897 VSS VSS nch l=0.04u w=0.8u
m1931 885 REFDIV[1] 69634 VSS nch l=0.04u w=0.8u
m1932 69637 930 886 VSS nch l=0.04u w=0.8u
m1933 VSS 485 69635 VSS nch l=0.04u w=0.8u
m1934 899 900 VSS VSS nch l=0.04u w=0.8u
m1935 901 902 VSS VSS nch l=0.04u w=0.8u
m1936 529 862 891 VSS nch l=0.04u w=0.4u
m1937 531 864 770 VSS nch l=0.04u w=0.4u
m1938 532 865 892 VSS nch l=0.04u w=0.4u
m1939 534 867 894 VSS nch l=0.04u w=0.4u
m1940 535 868 733 VSS nch l=0.04u w=0.4u
m1941 537 870 734 VSS nch l=0.04u w=0.4u
m1942 539 872 704 VSS nch l=0.04u w=0.4u
m1943 540 873 819 VSS nch l=0.04u w=0.4u
m1944 542 875 633 VSS nch l=0.04u w=0.4u
m1945 543 876 758 VSS nch l=0.04u w=0.4u
m1946 544 877 739 VSS nch l=0.04u w=0.4u
m1947 546 879 634 VSS nch l=0.04u w=0.4u
m1948 547 880 756 VSS nch l=0.04u w=0.4u
m1949 769 919 863 VSS nch l=0.04u w=0.4u
m1950 893 920 866 VSS nch l=0.04u w=0.4u
m1951 895 921 869 VSS nch l=0.04u w=0.4u
m1952 896 922 871 VSS nch l=0.04u w=0.4u
m1953 471 923 874 VSS nch l=0.04u w=0.4u
m1954 472 924 878 VSS nch l=0.04u w=0.4u
m1955 69639 858 VSS VSS nch l=0.04u w=0.8u
m1956 VSS 668 VSS VSS nch l=0.26u w=0.8u
m1957 VSS 671 VSS VSS nch l=0.26u w=0.8u
m1958 912 859 VSS VSS nch l=0.04u w=0.4u
m1959 913 860 VSS VSS nch l=0.04u w=0.4u
m1960 VSS 744 VSS VSS nch l=0.26u w=0.8u
m1961 914 4328 881 VSS nch l=0.04u w=0.4u
m1962 915 4328 882 VSS nch l=0.04u w=0.4u
m1963 916 4328 883 VSS nch l=0.04u w=0.4u
m1964 917 4328 884 VSS nch l=0.04u w=0.4u
m1965 VSS 2648 69637 VSS nch l=0.04u w=0.8u
m1966 VSS 909 909 VSS nch l=0.04u w=0.8u
m1967 919 863 769 VSS nch l=0.04u w=0.4u
m1968 920 866 893 VSS nch l=0.04u w=0.4u
m1969 921 869 895 VSS nch l=0.04u w=0.4u
m1970 922 871 896 VSS nch l=0.04u w=0.4u
m1971 923 874 471 VSS nch l=0.04u w=0.4u
m1972 924 878 472 VSS nch l=0.04u w=0.4u
m1973 911 817 69639 VSS nch l=0.04u w=0.8u
m1974 926 925 VSS VSS nch l=0.04u w=0.8u
m1975 927 928 VSS VSS nch l=0.04u w=0.8u
m1976 69664 806 914 VSS nch l=0.04u w=0.12u
m1977 69665 807 915 VSS nch l=0.04u w=0.12u
m1978 69666 808 916 VSS nch l=0.04u w=0.12u
m1979 69667 809 917 VSS nch l=0.04u w=0.12u
m1980 69668 853 VSS VSS nch l=0.04u w=0.8u
m1981 VSS 944 918 VSS nch l=0.04u w=0.4u
m1982 69671 1001 VSS VSS nch l=0.04u w=0.8u
m1983 VSS 903 919 VSS nch l=0.04u w=0.4u
m1984 69672 962 VSS VSS nch l=0.04u w=0.8u
m1985 VSS 904 920 VSS nch l=0.04u w=0.4u
m1986 VSS 905 921 VSS nch l=0.04u w=0.4u
m1987 VSS 906 922 VSS nch l=0.04u w=0.4u
m1988 VSS 907 923 VSS nch l=0.04u w=0.4u
m1989 VSS 908 924 VSS nch l=0.04u w=0.4u
m1990 VSS 744 VSS VSS nch l=0.26u w=0.8u
m1991 942 4328 VSS VSS nch l=0.04u w=0.4u
m1992 943 4328 VSS VSS nch l=0.04u w=0.4u
m1993 VSS 960 69664 VSS nch l=0.04u w=0.12u
m1994 VSS 737 69665 VSS nch l=0.04u w=0.12u
m1995 VSS 961 69666 VSS nch l=0.04u w=0.12u
m1996 VSS 740 69667 VSS nch l=0.04u w=0.12u
m1997 929 797 69668 VSS nch l=0.04u w=0.8u
m1998 VSS 966 930 VSS nch l=0.04u w=0.4u
m1999 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2000 931 979 69671 VSS nch l=0.04u w=0.8u
m2001 932 294 69672 VSS nch l=0.04u w=0.8u
m2002 VSS 933 933 VSS nch l=0.04u w=0.8u
m2003 69675 1041 VSS VSS nch l=0.04u w=0.8u
m2004 69676 1028 VSS VSS nch l=0.04u w=0.8u
m2005 69677 139 VSS VSS nch l=0.04u w=0.8u
m2006 69678 1042 VSS VSS nch l=0.04u w=0.8u
m2007 69679 2616 VSS VSS nch l=0.04u w=0.8u
m2008 69680 2616 VSS VSS nch l=0.04u w=0.8u
m2009 VSS 935 935 VSS nch l=0.04u w=0.8u
m2010 69681 1043 VSS VSS nch l=0.04u w=0.8u
m2011 69682 FRAC[3] VSS VSS nch l=0.04u w=0.8u
m2012 VSS 995 937 VSS nch l=0.04u w=0.4u
m2013 69683 1029 VSS VSS nch l=0.04u w=0.8u
m2014 69684 1045 VSS VSS nch l=0.04u w=0.8u
m2015 69685 998 VSS VSS nch l=0.04u w=0.8u
m2016 69686 937 VSS VSS nch l=0.04u w=0.8u
m2017 69687 1043 VSS VSS nch l=0.04u w=0.8u
m2018 69688 FRAC[3] VSS VSS nch l=0.04u w=0.8u
m2019 69689 937 VSS VSS nch l=0.04u w=0.8u
m2020 VSS 939 939 VSS nch l=0.04u w=0.8u
m2021 VSS 940 940 VSS nch l=0.04u w=0.8u
m2022 960 914 VSS VSS nch l=0.04u w=0.4u
m2023 737 915 VSS VSS nch l=0.04u w=0.4u
m2024 961 916 VSS VSS nch l=0.04u w=0.4u
m2025 740 917 VSS VSS nch l=0.04u w=0.4u
m2026 69690 854 VSS VSS nch l=0.04u w=0.12u
m2027 69691 2194 944 VSS nch l=0.04u w=0.8u
m2028 945 1023 69675 VSS nch l=0.04u w=0.8u
m2029 69694 1114 571 VSS nch l=0.04u w=0.8u
m2030 946 1024 69676 VSS nch l=0.04u w=0.8u
m2031 947 1025 69677 VSS nch l=0.04u w=0.8u
m2032 69695 1117 574 VSS nch l=0.04u w=0.8u
m2033 948 1026 69678 VSS nch l=0.04u w=0.8u
m2034 949 1182 69679 VSS nch l=0.04u w=0.8u
m2035 950 1183 69680 VSS nch l=0.04u w=0.8u
m2036 951 1027 69681 VSS nch l=0.04u w=0.8u
m2037 69696 1120 577 VSS nch l=0.04u w=0.8u
m2038 952 1028 69682 VSS nch l=0.04u w=0.8u
m2039 69697 1122 579 VSS nch l=0.04u w=0.8u
m2040 953 131 69683 VSS nch l=0.04u w=0.8u
m2041 954 1029 69684 VSS nch l=0.04u w=0.8u
m2042 69698 1125 582 VSS nch l=0.04u w=0.8u
m2043 955 1030 69685 VSS nch l=0.04u w=0.8u
m2044 956 999 69686 VSS nch l=0.04u w=0.8u
m2045 957 1031 69687 VSS nch l=0.04u w=0.8u
m2046 69699 1129 586 VSS nch l=0.04u w=0.8u
m2047 958 1032 69688 VSS nch l=0.04u w=0.8u
m2048 959 FBDIV[3] 69689 VSS nch l=0.04u w=0.8u
m2049 VSS 744 VSS VSS nch l=0.26u w=0.8u
m2050 963 942 912 VSS nch l=0.04u w=0.4u
m2051 964 943 913 VSS nch l=0.04u w=0.4u
m2052 966 1112 69690 VSS nch l=0.04u w=0.12u
m2053 69701 929 VSS VSS nch l=0.04u w=0.8u
m2054 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2055 69702 1653 69691 VSS nch l=0.04u w=0.8u
m2056 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2057 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2058 967 979 VSS VSS nch l=0.04u w=0.4u
m2059 VSS 1004 69694 VSS nch l=0.04u w=0.8u
m2060 968 294 VSS VSS nch l=0.04u w=0.4u
m2061 VSS 1007 69695 VSS nch l=0.04u w=0.8u
m2062 VSS 1010 69696 VSS nch l=0.04u w=0.8u
m2063 VSS 1013 69697 VSS nch l=0.04u w=0.8u
m2064 VSS 1016 69698 VSS nch l=0.04u w=0.8u
m2065 VSS 1020 69699 VSS nch l=0.04u w=0.8u
m2066 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2067 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2068 969 4328 VSS VSS nch l=0.04u w=0.4u
m2069 970 971 VSS VSS nch l=0.04u w=0.8u
m2070 VSS 2465 962 VSS nch l=0.04u w=0.4u
m2071 69705 4328 963 VSS nch l=0.04u w=0.12u
m2072 69706 4328 964 VSS nch l=0.04u w=0.12u
m2073 972 4328 VSS VSS nch l=0.04u w=0.4u
m2074 973 4328 VSS VSS nch l=0.04u w=0.4u
m2075 974 4328 VSS VSS nch l=0.04u w=0.4u
m2076 975 4328 VSS VSS nch l=0.04u w=0.4u
m2077 976 1152 966 VSS nch l=0.04u w=0.4u
m2078 965 885 69701 VSS nch l=0.04u w=0.8u
m2079 VSS 1061 69702 VSS nch l=0.04u w=0.8u
m2080 977 1001 967 VSS nch l=0.04u w=0.4u
m2081 978 962 968 VSS nch l=0.04u w=0.4u
m2082 980 1023 VSS VSS nch l=0.04u w=0.4u
m2083 981 1024 VSS VSS nch l=0.04u w=0.4u
m2084 982 1025 VSS VSS nch l=0.04u w=0.4u
m2085 983 1026 VSS VSS nch l=0.04u w=0.4u
m2086 984 949 VSS VSS nch l=0.04u w=0.4u
m2087 985 950 VSS VSS nch l=0.04u w=0.4u
m2088 986 1027 VSS VSS nch l=0.04u w=0.4u
m2089 987 1028 VSS VSS nch l=0.04u w=0.4u
m2090 988 131 VSS VSS nch l=0.04u w=0.4u
m2091 989 1029 VSS VSS nch l=0.04u w=0.4u
m2092 990 1030 VSS VSS nch l=0.04u w=0.4u
m2093 991 999 VSS VSS nch l=0.04u w=0.4u
m2094 992 1031 VSS VSS nch l=0.04u w=0.4u
m2095 993 1032 VSS VSS nch l=0.04u w=0.4u
m2096 994 FBDIV[3] VSS VSS nch l=0.04u w=0.4u
m2097 VSS 1035 69705 VSS nch l=0.04u w=0.12u
m2098 VSS 1036 69706 VSS nch l=0.04u w=0.12u
m2099 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2100 69711 885 965 VSS nch l=0.04u w=0.8u
m2101 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2102 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2103 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2104 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2105 1001 967 977 VSS nch l=0.04u w=0.4u
m2106 962 968 978 VSS nch l=0.04u w=0.4u
m2107 1003 1041 980 VSS nch l=0.04u w=0.4u
m2108 69712 863 VSS VSS nch l=0.04u w=0.8u
m2109 1005 1028 981 VSS nch l=0.04u w=0.4u
m2110 1006 139 982 VSS nch l=0.04u w=0.4u
m2111 69713 866 VSS VSS nch l=0.04u w=0.8u
m2112 1008 1042 983 VSS nch l=0.04u w=0.4u
m2113 1009 1043 986 VSS nch l=0.04u w=0.4u
m2114 69714 869 VSS VSS nch l=0.04u w=0.8u
m2115 1011 FRAC[3] 987 VSS nch l=0.04u w=0.4u
m2116 69715 871 VSS VSS nch l=0.04u w=0.8u
m2117 1014 1029 988 VSS nch l=0.04u w=0.4u
m2118 1015 1045 989 VSS nch l=0.04u w=0.4u
m2119 69716 874 VSS VSS nch l=0.04u w=0.8u
m2120 1017 998 990 VSS nch l=0.04u w=0.4u
m2121 1018 937 991 VSS nch l=0.04u w=0.4u
m2122 1019 1043 992 VSS nch l=0.04u w=0.4u
m2123 69717 878 VSS VSS nch l=0.04u w=0.8u
m2124 1021 FRAC[3] 993 VSS nch l=0.04u w=0.4u
m2125 1022 937 994 VSS nch l=0.04u w=0.4u
m2126 1012 969 995 VSS nch l=0.04u w=0.4u
m2127 1035 963 VSS VSS nch l=0.04u w=0.4u
m2128 1036 964 VSS VSS nch l=0.04u w=0.4u
m2129 1037 972 996 VSS nch l=0.04u w=0.4u
m2130 1038 973 997 VSS nch l=0.04u w=0.4u
m2131 1039 974 998 VSS nch l=0.04u w=0.4u
m2132 1040 975 999 VSS nch l=0.04u w=0.4u
m2133 VSS 929 69711 VSS nch l=0.04u w=0.8u
m2134 69721 1085 976 VSS nch l=0.04u w=0.8u
m2135 VSS 1240 1000 VSS nch l=0.04u w=0.4u
m2136 1041 980 1003 VSS nch l=0.04u w=0.4u
m2137 1004 903 69712 VSS nch l=0.04u w=0.8u
m2138 1028 981 1005 VSS nch l=0.04u w=0.4u
m2139 139 982 1006 VSS nch l=0.04u w=0.4u
m2140 1007 904 69713 VSS nch l=0.04u w=0.8u
m2141 1042 983 1008 VSS nch l=0.04u w=0.4u
m2142 1043 986 1009 VSS nch l=0.04u w=0.4u
m2143 1010 905 69714 VSS nch l=0.04u w=0.8u
m2144 FRAC[3] 987 1011 VSS nch l=0.04u w=0.4u
m2145 1013 906 69715 VSS nch l=0.04u w=0.8u
m2146 1029 988 1014 VSS nch l=0.04u w=0.4u
m2147 1045 989 1015 VSS nch l=0.04u w=0.4u
m2148 1016 907 69716 VSS nch l=0.04u w=0.8u
m2149 998 990 1017 VSS nch l=0.04u w=0.4u
m2150 937 991 1018 VSS nch l=0.04u w=0.4u
m2151 1043 992 1019 VSS nch l=0.04u w=0.4u
m2152 1020 908 69717 VSS nch l=0.04u w=0.8u
m2153 FRAC[3] 993 1021 VSS nch l=0.04u w=0.4u
m2154 937 994 1022 VSS nch l=0.04u w=0.4u
m2155 1046 1055 VSS VSS nch l=0.04u w=0.4u
m2156 1047 4328 VSS VSS nch l=0.04u w=0.4u
m2157 1048 4328 VSS VSS nch l=0.04u w=0.4u
m2158 1049 4328 VSS VSS nch l=0.04u w=0.4u
m2159 1050 4328 VSS VSS nch l=0.04u w=0.4u
m2160 69722 4328 1012 VSS nch l=0.04u w=0.12u
m2161 VSS 1080 1034 VSS nch l=0.04u w=0.4u
m2162 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2163 69728 4328 1037 VSS nch l=0.04u w=0.12u
m2164 69729 4328 1038 VSS nch l=0.04u w=0.12u
m2165 69730 4328 1039 VSS nch l=0.04u w=0.12u
m2166 69731 4328 1040 VSS nch l=0.04u w=0.12u
m2167 VSS 2648 69721 VSS nch l=0.04u w=0.8u
m2168 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2169 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2170 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2171 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2172 1051 1034 1046 VSS nch l=0.04u w=0.4u
m2173 VSS 1066 69722 VSS nch l=0.04u w=0.12u
m2174 69732 1034 VSS VSS nch l=0.04u w=0.12u
m2175 1058 4328 1035 VSS nch l=0.04u w=0.4u
m2176 1059 4328 1036 VSS nch l=0.04u w=0.4u
m2177 VSS 1081 69728 VSS nch l=0.04u w=0.12u
m2178 VSS 1082 69729 VSS nch l=0.04u w=0.12u
m2179 VSS 1083 69730 VSS nch l=0.04u w=0.12u
m2180 VSS 1084 69731 VSS nch l=0.04u w=0.12u
m2181 69752 976 VSS VSS nch l=0.04u w=0.24u
m2182 1060 76 VSS VSS nch l=0.04u w=0.4u
m2183 1061 1090 VSS VSS nch l=0.04u w=0.4u
m2184 1034 1046 1051 VSS nch l=0.04u w=0.4u
m2185 69755 977 1052 VSS nch l=0.04u w=0.8u
m2186 69756 978 1053 VSS nch l=0.04u w=0.8u
m2187 1066 1012 VSS VSS nch l=0.04u w=0.4u
m2188 1062 1047 1056 VSS nch l=0.04u w=0.4u
m2189 1063 1048 1057 VSS nch l=0.04u w=0.4u
m2190 1064 1049 984 VSS nch l=0.04u w=0.4u
m2191 1065 1050 985 VSS nch l=0.04u w=0.4u
m2192 1080 1176 69732 VSS nch l=0.04u w=0.12u
m2193 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2194 69757 942 1058 VSS nch l=0.04u w=0.12u
m2195 69758 943 1059 VSS nch l=0.04u w=0.12u
m2196 1081 1037 VSS VSS nch l=0.04u w=0.4u
m2197 1082 1038 VSS VSS nch l=0.04u w=0.4u
m2198 1083 1039 VSS VSS nch l=0.04u w=0.4u
m2199 1084 1040 VSS VSS nch l=0.04u w=0.4u
m2200 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2201 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2202 1085 1152 69752 VSS nch l=0.04u w=0.24u
m2203 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2204 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2205 VSS 1090 1061 VSS nch l=0.04u w=0.4u
m2206 VSS 811 69755 VSS nch l=0.04u w=0.8u
m2207 VSS 814 69756 VSS nch l=0.04u w=0.8u
m2208 69759 4328 1062 VSS nch l=0.04u w=0.12u
m2209 69760 4328 1063 VSS nch l=0.04u w=0.12u
m2210 69761 1003 1067 VSS nch l=0.04u w=0.8u
m2211 903 1092 569 VSS nch l=0.04u w=0.4u
m2212 69762 1005 1068 VSS nch l=0.04u w=0.8u
m2213 69763 1006 1069 VSS nch l=0.04u w=0.8u
m2214 904 1093 139 VSS nch l=0.04u w=0.4u
m2215 69764 1008 1070 VSS nch l=0.04u w=0.8u
m2216 69765 4328 1064 VSS nch l=0.04u w=0.12u
m2217 69766 4328 1065 VSS nch l=0.04u w=0.12u
m2218 69767 1009 1071 VSS nch l=0.04u w=0.8u
m2219 905 1094 FRAC[21] VSS nch l=0.04u w=0.4u
m2220 69768 1011 1072 VSS nch l=0.04u w=0.8u
m2221 906 1095 589 VSS nch l=0.04u w=0.4u
m2222 69769 1014 1073 VSS nch l=0.04u w=0.8u
m2223 69770 1015 1074 VSS nch l=0.04u w=0.8u
m2224 907 1096 472 VSS nch l=0.04u w=0.4u
m2225 69771 1017 1075 VSS nch l=0.04u w=0.8u
m2226 69772 1018 1076 VSS nch l=0.04u w=0.8u
m2227 69773 1019 1077 VSS nch l=0.04u w=0.8u
m2228 908 1097 FRAC[21] VSS nch l=0.04u w=0.4u
m2229 69774 1021 1078 VSS nch l=0.04u w=0.8u
m2230 69775 1022 1079 VSS nch l=0.04u w=0.8u
m2231 1087 1593 1080 VSS nch l=0.04u w=0.4u
m2232 1088 155 VSS VSS nch l=0.04u w=0.4u
m2233 VSS 1098 69757 VSS nch l=0.04u w=0.12u
m2234 VSS 1099 69758 VSS nch l=0.04u w=0.12u
m2235 886 1112 1085 VSS nch l=0.04u w=0.4u
m2236 1089 1060 965 VSS nch l=0.04u w=0.4u
m2237 VSS 1105 69759 VSS nch l=0.04u w=0.12u
m2238 VSS 1106 69760 VSS nch l=0.04u w=0.12u
m2239 VSS 822 69761 VSS nch l=0.04u w=0.8u
m2240 1092 569 903 VSS nch l=0.04u w=0.4u
m2241 VSS 824 69762 VSS nch l=0.04u w=0.8u
m2242 VSS 825 69763 VSS nch l=0.04u w=0.8u
m2243 1093 139 904 VSS nch l=0.04u w=0.4u
m2244 VSS 827 69764 VSS nch l=0.04u w=0.8u
m2245 VSS 1108 69765 VSS nch l=0.04u w=0.12u
m2246 VSS 1109 69766 VSS nch l=0.04u w=0.12u
m2247 VSS 828 69767 VSS nch l=0.04u w=0.8u
m2248 1094 FRAC[21] 905 VSS nch l=0.04u w=0.4u
m2249 VSS 830 69768 VSS nch l=0.04u w=0.8u
m2250 1091 4328 1066 VSS nch l=0.04u w=0.4u
m2251 1095 589 906 VSS nch l=0.04u w=0.4u
m2252 VSS 832 69769 VSS nch l=0.04u w=0.8u
m2253 VSS 833 69770 VSS nch l=0.04u w=0.8u
m2254 1096 472 907 VSS nch l=0.04u w=0.4u
m2255 VSS 835 69771 VSS nch l=0.04u w=0.8u
m2256 VSS 836 69772 VSS nch l=0.04u w=0.8u
m2257 VSS 837 69773 VSS nch l=0.04u w=0.8u
m2258 1097 FRAC[21] 908 VSS nch l=0.04u w=0.4u
m2259 VSS 839 69774 VSS nch l=0.04u w=0.8u
m2260 VSS 840 69775 VSS nch l=0.04u w=0.8u
m2261 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2262 1098 1058 VSS VSS nch l=0.04u w=0.4u
m2263 1099 1059 VSS VSS nch l=0.04u w=0.4u
m2264 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2265 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2266 1100 4328 1081 VSS nch l=0.04u w=0.4u
m2267 1101 4328 1082 VSS nch l=0.04u w=0.4u
m2268 1102 4328 1083 VSS nch l=0.04u w=0.4u
m2269 1103 4328 1084 VSS nch l=0.04u w=0.4u
m2270 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2271 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2272 69779 76 1089 VSS nch l=0.04u w=0.12u
m2273 VSS 1137 1090 VSS nch l=0.04u w=0.4u
m2274 69780 1052 VSS VSS nch l=0.04u w=0.8u
m2275 1105 1062 VSS VSS nch l=0.04u w=0.4u
m2276 1106 1063 VSS VSS nch l=0.04u w=0.4u
m2277 VSS 888 1092 VSS nch l=0.04u w=0.4u
m2278 69781 1053 VSS VSS nch l=0.04u w=0.8u
m2279 VSS 895 1093 VSS nch l=0.04u w=0.4u
m2280 1108 1064 VSS VSS nch l=0.04u w=0.4u
m2281 1109 1065 VSS VSS nch l=0.04u w=0.4u
m2282 VSS 398 1094 VSS nch l=0.04u w=0.4u
m2283 69782 969 1091 VSS nch l=0.04u w=0.12u
m2284 VSS 1086 1095 VSS nch l=0.04u w=0.4u
m2285 VSS 589 1096 VSS nch l=0.04u w=0.4u
m2286 VSS 590 1097 VSS nch l=0.04u w=0.4u
m2287 1110 PD VSS VSS nch l=0.04u w=0.4u
m2288 VSS 1143 1087 VSS nch l=0.04u w=0.4u
m2289 69783 155 VSS VSS nch l=0.04u w=0.8u
m2290 69784 972 1100 VSS nch l=0.04u w=0.12u
m2291 69785 973 1101 VSS nch l=0.04u w=0.12u
m2292 69786 974 1102 VSS nch l=0.04u w=0.12u
m2293 69787 975 1103 VSS nch l=0.04u w=0.12u
m2294 1112 1152 VSS VSS nch l=0.04u w=0.4u
m2295 VSS 1135 69779 VSS nch l=0.04u w=0.12u
m2296 69788 1090 VSS VSS nch l=0.04u w=0.12u
m2297 1104 931 69780 VSS nch l=0.04u w=0.8u
m2298 1107 932 69781 VSS nch l=0.04u w=0.8u
m2299 VSS 1142 69782 VSS nch l=0.04u w=0.12u
m2300 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2301 69791 1067 VSS VSS nch l=0.04u w=0.8u
m2302 69792 1068 VSS VSS nch l=0.04u w=0.8u
m2303 69793 1069 VSS VSS nch l=0.04u w=0.8u
m2304 69794 1070 VSS VSS nch l=0.04u w=0.8u
m2305 69795 1071 VSS VSS nch l=0.04u w=0.8u
m2306 69796 1072 VSS VSS nch l=0.04u w=0.8u
m2307 69797 1073 VSS VSS nch l=0.04u w=0.8u
m2308 69798 1074 VSS VSS nch l=0.04u w=0.8u
m2309 69799 1075 VSS VSS nch l=0.04u w=0.8u
m2310 69800 1076 VSS VSS nch l=0.04u w=0.8u
m2311 69801 1077 VSS VSS nch l=0.04u w=0.8u
m2312 69802 1078 VSS VSS nch l=0.04u w=0.8u
m2313 69803 1079 VSS VSS nch l=0.04u w=0.8u
m2314 69804 1087 VSS VSS nch l=0.04u w=0.12u
m2315 1111 FBDIV[3] 69783 VSS nch l=0.04u w=0.8u
m2316 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2317 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2318 1133 1146 VSS VSS nch l=0.04u w=0.4u
m2319 1134 70 VSS VSS nch l=0.04u w=0.4u
m2320 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2321 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2322 VSS 1030 69784 VSS nch l=0.04u w=0.12u
m2323 VSS 1029 69785 VSS nch l=0.04u w=0.12u
m2324 VSS 1032 69786 VSS nch l=0.04u w=0.12u
m2325 VSS 1031 69787 VSS nch l=0.04u w=0.12u
m2326 1135 1089 VSS VSS nch l=0.04u w=0.4u
m2327 1137 1241 69788 VSS nch l=0.04u w=0.12u
m2328 1142 1091 VSS VSS nch l=0.04u w=0.4u
m2329 1138 4328 1105 VSS nch l=0.04u w=0.4u
m2330 1139 4328 1106 VSS nch l=0.04u w=0.4u
m2331 1113 945 69791 VSS nch l=0.04u w=0.8u
m2332 69805 888 1114 VSS nch l=0.04u w=0.8u
m2333 1115 946 69792 VSS nch l=0.04u w=0.8u
m2334 1116 947 69793 VSS nch l=0.04u w=0.8u
m2335 69806 895 1117 VSS nch l=0.04u w=0.8u
m2336 1118 948 69794 VSS nch l=0.04u w=0.8u
m2337 1140 4328 1108 VSS nch l=0.04u w=0.4u
m2338 1141 4328 1109 VSS nch l=0.04u w=0.4u
m2339 1119 951 69795 VSS nch l=0.04u w=0.8u
m2340 69807 398 1120 VSS nch l=0.04u w=0.8u
m2341 1121 952 69796 VSS nch l=0.04u w=0.8u
m2342 69808 1086 1122 VSS nch l=0.04u w=0.8u
m2343 1123 953 69797 VSS nch l=0.04u w=0.8u
m2344 1124 954 69798 VSS nch l=0.04u w=0.8u
m2345 69809 589 1125 VSS nch l=0.04u w=0.8u
m2346 1126 955 69799 VSS nch l=0.04u w=0.8u
m2347 1127 956 69800 VSS nch l=0.04u w=0.8u
m2348 1128 957 69801 VSS nch l=0.04u w=0.8u
m2349 69810 590 1129 VSS nch l=0.04u w=0.8u
m2350 1130 958 69802 VSS nch l=0.04u w=0.8u
m2351 1131 959 69803 VSS nch l=0.04u w=0.8u
m2352 1143 1593 69804 VSS nch l=0.04u w=0.12u
m2353 VSS 1372 1132 VSS nch l=0.04u w=0.4u
m2354 1144 1098 1133 VSS nch l=0.04u w=0.4u
m2355 1145 1099 1134 VSS nch l=0.04u w=0.4u
m2356 1030 1100 VSS VSS nch l=0.04u w=0.4u
m2357 1029 1101 VSS VSS nch l=0.04u w=0.4u
m2358 1032 1102 VSS VSS nch l=0.04u w=0.4u
m2359 1031 1103 VSS VSS nch l=0.04u w=0.4u
m2360 VSS 1152 1136 VSS nch l=0.04u w=0.4u
m2361 1147 76 1137 VSS nch l=0.04u w=0.4u
m2362 VSS 910 VSS VSS nch l=0.26u w=0.8u
m2363 1148 977 VSS VSS nch l=0.04u w=0.4u
m2364 69813 1047 1138 VSS nch l=0.04u w=0.12u
m2365 69814 1048 1139 VSS nch l=0.04u w=0.12u
m2366 VSS 569 69805 VSS nch l=0.04u w=0.8u
m2367 1149 978 VSS VSS nch l=0.04u w=0.4u
m2368 VSS 139 69806 VSS nch l=0.04u w=0.8u
m2369 69815 1049 1140 VSS nch l=0.04u w=0.12u
m2370 69816 1050 1141 VSS nch l=0.04u w=0.12u
m2371 VSS FRAC[21] 69807 VSS nch l=0.04u w=0.8u
m2372 VSS 589 69808 VSS nch l=0.04u w=0.8u
m2373 VSS 472 69809 VSS nch l=0.04u w=0.8u
m2374 VSS FRAC[21] 69810 VSS nch l=0.04u w=0.8u
m2375 1055 1176 1143 VSS nch l=0.04u w=0.4u
m2376 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2377 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2378 69817 1088 VSS VSS nch l=0.04u w=0.8u
m2379 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2380 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2381 1098 1133 1144 VSS nch l=0.04u w=0.4u
m2382 1099 1134 1145 VSS nch l=0.04u w=0.4u
m2383 1151 76 1135 VSS nch l=0.04u w=0.4u
m2384 1153 1154 VSS VSS nch l=0.04u w=0.8u
m2385 1155 811 1148 VSS nch l=0.04u w=0.4u
m2386 VSS 1179 69813 VSS nch l=0.04u w=0.12u
m2387 VSS 1024 69814 VSS nch l=0.04u w=0.12u
m2388 474 814 1149 VSS nch l=0.04u w=0.4u
m2389 VSS 94 69815 VSS nch l=0.04u w=0.12u
m2390 VSS 1028 69816 VSS nch l=0.04u w=0.12u
m2391 1156 1156 VSS VSS nch l=0.04u w=0.8u
m2392 1158 1003 VSS VSS nch l=0.04u w=0.4u
m2393 1160 1005 VSS VSS nch l=0.04u w=0.4u
m2394 1161 1006 VSS VSS nch l=0.04u w=0.4u
m2395 1163 1008 VSS VSS nch l=0.04u w=0.4u
m2396 1164 1009 VSS VSS nch l=0.04u w=0.4u
m2397 1166 1011 VSS VSS nch l=0.04u w=0.4u
m2398 1167 1014 VSS VSS nch l=0.04u w=0.4u
m2399 1168 1015 VSS VSS nch l=0.04u w=0.4u
m2400 1170 1017 VSS VSS nch l=0.04u w=0.4u
m2401 1171 1018 VSS VSS nch l=0.04u w=0.4u
m2402 1172 1019 VSS VSS nch l=0.04u w=0.4u
m2403 1174 1021 VSS VSS nch l=0.04u w=0.4u
m2404 1175 1022 VSS VSS nch l=0.04u w=0.4u
m2405 1157 1132 1051 VSS nch l=0.04u w=0.4u
m2406 1150 1142 69817 VSS nch l=0.04u w=0.8u
m2407 69828 1060 1151 VSS nch l=0.04u w=0.12u
m2408 69829 1201 1152 VSS nch l=0.04u w=0.8u
m2409 VSS 1202 1147 VSS nch l=0.04u w=0.4u
m2410 811 1148 1155 VSS nch l=0.04u w=0.4u
m2411 1179 1138 VSS VSS nch l=0.04u w=0.4u
m2412 1024 1139 VSS VSS nch l=0.04u w=0.4u
m2413 VSS 934 VSS VSS nch l=0.26u w=0.8u
m2414 814 1149 474 VSS nch l=0.04u w=0.4u
m2415 94 1140 VSS VSS nch l=0.04u w=0.4u
m2416 1028 1141 VSS VSS nch l=0.04u w=0.4u
m2417 VSS 936 VSS VSS nch l=0.26u w=0.8u
m2418 1180 822 1158 VSS nch l=0.04u w=0.4u
m2419 1057 824 1160 VSS nch l=0.04u w=0.4u
m2420 1181 825 1161 VSS nch l=0.04u w=0.4u
m2421 1183 827 1163 VSS nch l=0.04u w=0.4u
m2422 1025 828 1164 VSS nch l=0.04u w=0.4u
m2423 1026 830 1166 VSS nch l=0.04u w=0.4u
m2424 995 832 1167 VSS nch l=0.04u w=0.4u
m2425 997 833 1168 VSS nch l=0.04u w=0.4u
m2426 996 835 1170 VSS nch l=0.04u w=0.4u
m2427 1045 836 1171 VSS nch l=0.04u w=0.4u
m2428 999 837 1172 VSS nch l=0.04u w=0.4u
m2429 998 839 1174 VSS nch l=0.04u w=0.4u
m2430 1043 840 1175 VSS nch l=0.04u w=0.4u
m2431 VSS 1593 1176 VSS nch l=0.04u w=0.4u
m2432 69834 1372 1157 VSS nch l=0.04u w=0.24u
m2433 VSS 938 VSS VSS nch l=0.26u w=0.8u
m2434 VSS 941 VSS VSS nch l=0.26u w=0.8u
m2435 VSS 810 69828 VSS nch l=0.04u w=0.12u
m2436 VSS 2648 69829 VSS nch l=0.04u w=0.8u
m2437 69835 1147 VSS VSS nch l=0.04u w=0.12u
m2438 VSS 1177 1177 VSS nch l=0.04u w=0.8u
m2439 1186 1187 VSS VSS nch l=0.04u w=0.8u
m2440 1188 1189 VSS VSS nch l=0.04u w=0.8u
m2441 822 1158 1180 VSS nch l=0.04u w=0.4u
m2442 824 1160 1057 VSS nch l=0.04u w=0.4u
m2443 825 1161 1181 VSS nch l=0.04u w=0.4u
m2444 827 1163 1183 VSS nch l=0.04u w=0.4u
m2445 828 1164 1025 VSS nch l=0.04u w=0.4u
m2446 830 1166 1026 VSS nch l=0.04u w=0.4u
m2447 832 1167 995 VSS nch l=0.04u w=0.4u
m2448 833 1168 997 VSS nch l=0.04u w=0.4u
m2449 835 1170 996 VSS nch l=0.04u w=0.4u
m2450 836 1171 1045 VSS nch l=0.04u w=0.4u
m2451 837 1172 999 VSS nch l=0.04u w=0.4u
m2452 839 1174 998 VSS nch l=0.04u w=0.4u
m2453 840 1175 1043 VSS nch l=0.04u w=0.4u
m2454 VSS 1204 69834 VSS nch l=0.04u w=0.24u
m2455 1197 1196 VSS VSS nch l=0.04u w=0.8u
m2456 1198 1199 VSS VSS nch l=0.04u w=0.8u
m2457 1056 1205 1159 VSS nch l=0.04u w=0.4u
m2458 1182 1206 1162 VSS nch l=0.04u w=0.4u
m2459 1184 1207 1165 VSS nch l=0.04u w=0.4u
m2460 1185 1208 131 VSS nch l=0.04u w=0.4u
m2461 818 1213 1169 VSS nch l=0.04u w=0.4u
m2462 820 1218 1173 VSS nch l=0.04u w=0.4u
m2463 69836 1150 VSS VSS nch l=0.04u w=0.8u
m2464 810 1151 VSS VSS nch l=0.04u w=0.4u
m2465 1202 76 69835 VSS nch l=0.04u w=0.12u
m2466 131 1203 VSS VSS nch l=0.04u w=0.8u
m2467 69843 1110 VSS VSS nch l=0.04u w=0.8u
m2468 1205 1159 1056 VSS nch l=0.04u w=0.4u
m2469 1206 1162 1182 VSS nch l=0.04u w=0.4u
m2470 1207 1165 1184 VSS nch l=0.04u w=0.4u
m2471 1208 131 1185 VSS nch l=0.04u w=0.4u
m2472 1213 1169 818 VSS nch l=0.04u w=0.4u
m2473 1218 1173 820 VSS nch l=0.04u w=0.4u
m2474 VSS 1257 1055 VSS nch l=0.04u w=0.4u
m2475 1200 1111 69836 VSS nch l=0.04u w=0.8u
m2476 1223 4328 VSS VSS nch l=0.04u w=0.4u
m2477 1224 4328 VSS VSS nch l=0.04u w=0.4u
m2478 VSS 1258 1201 VSS nch l=0.04u w=0.4u
m2479 1225 1241 1202 VSS nch l=0.04u w=0.4u
m2480 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2481 1204 1157 69843 VSS nch l=0.04u w=0.8u
m2482 1226 1104 VSS VSS nch l=0.04u w=0.4u
m2483 VSS 1190 1205 VSS nch l=0.04u w=0.4u
m2484 1227 1107 VSS VSS nch l=0.04u w=0.4u
m2485 VSS 1191 1206 VSS nch l=0.04u w=0.4u
m2486 VSS 1192 1207 VSS nch l=0.04u w=0.4u
m2487 VSS 1193 1208 VSS nch l=0.04u w=0.4u
m2488 VSS 1210 1210 VSS nch l=0.04u w=0.8u
m2489 VSS 1211 1211 VSS nch l=0.04u w=0.8u
m2490 VSS 1194 1213 VSS nch l=0.04u w=0.4u
m2491 VSS 1215 1215 VSS nch l=0.04u w=0.8u
m2492 VSS 1216 1216 VSS nch l=0.04u w=0.8u
m2493 VSS 1195 1218 VSS nch l=0.04u w=0.4u
m2494 69863 1055 VSS VSS nch l=0.04u w=0.12u
m2495 VSS 1220 1220 VSS nch l=0.04u w=0.8u
m2496 VSS 1221 1221 VSS nch l=0.04u w=0.8u
m2497 1240 810 VSS VSS nch l=0.04u w=0.4u
m2498 69865 1136 VSS VSS nch l=0.04u w=0.12u
m2499 1257 1315 69863 VSS nch l=0.04u w=0.12u
m2500 1242 1113 VSS VSS nch l=0.04u w=0.4u
m2501 1243 1115 VSS VSS nch l=0.04u w=0.4u
m2502 1244 1116 VSS VSS nch l=0.04u w=0.4u
m2503 1245 1118 VSS VSS nch l=0.04u w=0.4u
m2504 1246 1119 VSS VSS nch l=0.04u w=0.4u
m2505 1247 1121 VSS VSS nch l=0.04u w=0.4u
m2506 1250 1123 VSS VSS nch l=0.04u w=0.4u
m2507 1251 1124 VSS VSS nch l=0.04u w=0.4u
m2508 1252 1126 VSS VSS nch l=0.04u w=0.4u
m2509 1253 1127 VSS VSS nch l=0.04u w=0.4u
m2510 1254 1128 VSS VSS nch l=0.04u w=0.4u
m2511 1255 1130 VSS VSS nch l=0.04u w=0.4u
m2512 1256 1131 VSS VSS nch l=0.04u w=0.4u
m2513 1248 1223 1144 VSS nch l=0.04u w=0.4u
m2514 1249 1224 1145 VSS nch l=0.04u w=0.4u
m2515 VSS 1228 1228 VSS nch l=0.04u w=0.8u
m2516 VSS 1231 1231 VSS nch l=0.04u w=0.8u
m2517 VSS 1232 1232 VSS nch l=0.04u w=0.8u
m2518 VSS 1234 1234 VSS nch l=0.04u w=0.8u
m2519 VSS 1237 1237 VSS nch l=0.04u w=0.8u
m2520 VSS 1238 1238 VSS nch l=0.04u w=0.8u
m2521 VSS 810 1240 VSS nch l=0.04u w=0.4u
m2522 1258 1353 69865 VSS nch l=0.04u w=0.12u
m2523 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2524 VSS 76 1241 VSS nch l=0.04u w=0.4u
m2525 VSS 1209 VSS VSS nch l=0.26u w=0.8u
m2526 VSS 1212 VSS VSS nch l=0.26u w=0.8u
m2527 VSS 1214 VSS VSS nch l=0.26u w=0.8u
m2528 VSS 1217 VSS VSS nch l=0.26u w=0.8u
m2529 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2530 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2531 1260 1372 1257 VSS nch l=0.04u w=0.4u
m2532 1259 1372 1204 VSS nch l=0.04u w=0.4u
m2533 69868 89 VSS VSS nch l=0.04u w=0.8u
m2534 69869 1373 863 VSS nch l=0.04u w=0.8u
m2535 69870 90 VSS VSS nch l=0.04u w=0.8u
m2536 69871 1374 866 VSS nch l=0.04u w=0.8u
m2537 69872 1375 869 VSS nch l=0.04u w=0.8u
m2538 69873 1376 871 VSS nch l=0.04u w=0.8u
m2539 69874 1377 874 VSS nch l=0.04u w=0.8u
m2540 69875 1378 878 VSS nch l=0.04u w=0.8u
m2541 69876 4328 1248 VSS nch l=0.04u w=0.12u
m2542 69877 4328 1249 VSS nch l=0.04u w=0.12u
m2543 1266 1392 1258 VSS nch l=0.04u w=0.4u
m2544 69879 1132 1259 VSS nch l=0.04u w=0.12u
m2545 69880 393 69868 VSS nch l=0.04u w=0.8u
m2546 VSS 1284 69869 VSS nch l=0.04u w=0.8u
m2547 69881 394 69870 VSS nch l=0.04u w=0.8u
m2548 VSS 1285 69871 VSS nch l=0.04u w=0.8u
m2549 VSS 1286 69872 VSS nch l=0.04u w=0.8u
m2550 VSS 1287 69873 VSS nch l=0.04u w=0.8u
m2551 VSS 1288 69874 VSS nch l=0.04u w=0.8u
m2552 VSS 1289 69875 VSS nch l=0.04u w=0.8u
m2553 69882 111 VSS VSS nch l=0.04u w=0.8u
m2554 69883 112 VSS VSS nch l=0.04u w=0.8u
m2555 69884 113 VSS VSS nch l=0.04u w=0.8u
m2556 69885 114 VSS VSS nch l=0.04u w=0.8u
m2557 69886 115 VSS VSS nch l=0.04u w=0.8u
m2558 69887 116 VSS VSS nch l=0.04u w=0.8u
m2559 VSS 1281 69876 VSS nch l=0.04u w=0.12u
m2560 VSS 1282 69877 VSS nch l=0.04u w=0.12u
m2561 69888 118 VSS VSS nch l=0.04u w=0.8u
m2562 69889 119 VSS VSS nch l=0.04u w=0.8u
m2563 69890 120 VSS VSS nch l=0.04u w=0.8u
m2564 69891 121 VSS VSS nch l=0.04u w=0.8u
m2565 69892 122 VSS VSS nch l=0.04u w=0.8u
m2566 69893 123 VSS VSS nch l=0.04u w=0.8u
m2567 69894 124 VSS VSS nch l=0.04u w=0.8u
m2568 VSS 1265 1265 VSS nch l=0.04u w=0.8u
m2569 VSS 1229 VSS VSS nch l=0.26u w=0.8u
m2570 VSS 1230 VSS VSS nch l=0.26u w=0.8u
m2571 VSS 1233 VSS VSS nch l=0.26u w=0.8u
m2572 VSS 1235 VSS VSS nch l=0.26u w=0.8u
m2573 VSS 1236 VSS VSS nch l=0.26u w=0.8u
m2574 VSS 1239 VSS VSS nch l=0.26u w=0.8u
m2575 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2576 69895 1240 VSS VSS nch l=0.04u w=0.8u
m2577 69896 1314 VSS VSS nch l=0.04u w=0.8u
m2578 VSS 1209 VSS VSS nch l=0.26u w=0.8u
m2579 VSS 1212 VSS VSS nch l=0.26u w=0.8u
m2580 VSS 1214 VSS VSS nch l=0.26u w=0.8u
m2581 VSS 1217 VSS VSS nch l=0.26u w=0.8u
m2582 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2583 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2584 VSS 1335 69879 VSS nch l=0.04u w=0.12u
m2585 1261 686 69880 VSS nch l=0.04u w=0.8u
m2586 1262 687 69881 VSS nch l=0.04u w=0.8u
m2587 VSS 1294 1260 VSS nch l=0.04u w=0.4u
m2588 69898 417 69882 VSS nch l=0.04u w=0.8u
m2589 69899 419 69883 VSS nch l=0.04u w=0.8u
m2590 69900 420 69884 VSS nch l=0.04u w=0.8u
m2591 69901 422 69885 VSS nch l=0.04u w=0.8u
m2592 69902 423 69886 VSS nch l=0.04u w=0.8u
m2593 69903 425 69887 VSS nch l=0.04u w=0.8u
m2594 1281 1248 VSS VSS nch l=0.04u w=0.4u
m2595 1282 1249 VSS VSS nch l=0.04u w=0.4u
m2596 69904 428 69888 VSS nch l=0.04u w=0.8u
m2597 69905 429 69889 VSS nch l=0.04u w=0.8u
m2598 69906 431 69890 VSS nch l=0.04u w=0.8u
m2599 69907 432 69891 VSS nch l=0.04u w=0.8u
m2600 69908 433 69892 VSS nch l=0.04u w=0.8u
m2601 69909 435 69893 VSS nch l=0.04u w=0.8u
m2602 69910 436 69894 VSS nch l=0.04u w=0.8u
m2603 1280 683 69895 VSS nch l=0.04u w=0.8u
m2604 69911 1313 1266 VSS nch l=0.04u w=0.8u
m2605 1225 1354 69896 VSS nch l=0.04u w=0.8u
m2606 1283 1259 VSS VSS nch l=0.04u w=0.4u
m2607 69912 1260 VSS VSS nch l=0.04u w=0.12u
m2608 1267 711 69898 VSS nch l=0.04u w=0.8u
m2609 69913 1159 VSS VSS nch l=0.04u w=0.8u
m2610 1268 713 69899 VSS nch l=0.04u w=0.8u
m2611 1269 714 69900 VSS nch l=0.04u w=0.8u
m2612 69914 1162 VSS VSS nch l=0.04u w=0.8u
m2613 1270 716 69901 VSS nch l=0.04u w=0.8u
m2614 1271 717 69902 VSS nch l=0.04u w=0.8u
m2615 69915 1165 VSS VSS nch l=0.04u w=0.8u
m2616 1272 719 69903 VSS nch l=0.04u w=0.8u
m2617 69916 131 VSS VSS nch l=0.04u w=0.8u
m2618 1273 722 69904 VSS nch l=0.04u w=0.8u
m2619 1274 723 69905 VSS nch l=0.04u w=0.8u
m2620 69917 1169 VSS VSS nch l=0.04u w=0.8u
m2621 1275 725 69906 VSS nch l=0.04u w=0.8u
m2622 1276 726 69907 VSS nch l=0.04u w=0.8u
m2623 1277 727 69908 VSS nch l=0.04u w=0.8u
m2624 69918 1173 VSS VSS nch l=0.04u w=0.8u
m2625 1278 729 69909 VSS nch l=0.04u w=0.8u
m2626 1279 730 69910 VSS nch l=0.04u w=0.8u
m2627 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2628 VSS 1229 VSS VSS nch l=0.26u w=0.8u
m2629 VSS 1230 VSS VSS nch l=0.26u w=0.8u
m2630 VSS 1233 VSS VSS nch l=0.26u w=0.8u
m2631 VSS 1235 VSS VSS nch l=0.26u w=0.8u
m2632 VSS 1236 VSS VSS nch l=0.26u w=0.8u
m2633 VSS 1239 VSS VSS nch l=0.26u w=0.8u
m2634 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2635 VSS 2648 69911 VSS nch l=0.04u w=0.8u
m2636 VSS 1209 VSS VSS nch l=0.26u w=0.8u
m2637 VSS 1212 VSS VSS nch l=0.26u w=0.8u
m2638 VSS 1214 VSS VSS nch l=0.26u w=0.8u
m2639 VSS 1217 VSS VSS nch l=0.26u w=0.8u
m2640 69919 1354 1225 VSS nch l=0.04u w=0.8u
m2641 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2642 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2643 1294 1372 69912 VSS nch l=0.04u w=0.12u
m2644 1290 1261 VSS VSS nch l=0.04u w=0.4u
m2645 1284 1190 69913 VSS nch l=0.04u w=0.8u
m2646 1291 1262 VSS VSS nch l=0.04u w=0.4u
m2647 1285 1191 69914 VSS nch l=0.04u w=0.8u
m2648 1286 1192 69915 VSS nch l=0.04u w=0.8u
m2649 1287 1193 69916 VSS nch l=0.04u w=0.8u
m2650 1288 1194 69917 VSS nch l=0.04u w=0.8u
m2651 1289 1195 69918 VSS nch l=0.04u w=0.8u
m2652 1292 4328 1281 VSS nch l=0.04u w=0.4u
m2653 1293 4328 1282 VSS nch l=0.04u w=0.4u
m2654 69921 1266 VSS VSS nch l=0.04u w=0.24u
m2655 1295 1280 VSS VSS nch l=0.04u w=0.4u
m2656 VSS 1314 69919 VSS nch l=0.04u w=0.8u
m2657 1296 1315 1294 VSS nch l=0.04u w=0.4u
m2658 69923 1110 VSS VSS nch l=0.04u w=0.8u
m2659 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2660 VSS 1229 VSS VSS nch l=0.26u w=0.8u
m2661 VSS 1230 VSS VSS nch l=0.26u w=0.8u
m2662 VSS 1233 VSS VSS nch l=0.26u w=0.8u
m2663 VSS 1235 VSS VSS nch l=0.26u w=0.8u
m2664 VSS 1236 VSS VSS nch l=0.26u w=0.8u
m2665 VSS 1239 VSS VSS nch l=0.26u w=0.8u
m2666 1298 1267 VSS VSS nch l=0.04u w=0.4u
m2667 1299 1268 VSS VSS nch l=0.04u w=0.4u
m2668 1300 1269 VSS VSS nch l=0.04u w=0.4u
m2669 1301 1270 VSS VSS nch l=0.04u w=0.4u
m2670 1302 1271 VSS VSS nch l=0.04u w=0.4u
m2671 1304 1272 VSS VSS nch l=0.04u w=0.4u
m2672 69924 1223 1292 VSS nch l=0.04u w=0.12u
m2673 69925 1224 1293 VSS nch l=0.04u w=0.12u
m2674 1305 1273 VSS VSS nch l=0.04u w=0.4u
m2675 1306 1274 VSS VSS nch l=0.04u w=0.4u
m2676 1307 1275 VSS VSS nch l=0.04u w=0.4u
m2677 1308 1276 VSS VSS nch l=0.04u w=0.4u
m2678 1309 1277 VSS VSS nch l=0.04u w=0.4u
m2679 1310 1278 VSS VSS nch l=0.04u w=0.4u
m2680 1311 1279 VSS VSS nch l=0.04u w=0.4u
m2681 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2682 1313 1392 69921 VSS nch l=0.04u w=0.24u
m2683 VSS 1209 VSS VSS nch l=0.26u w=0.8u
m2684 VSS 1212 VSS VSS nch l=0.26u w=0.8u
m2685 VSS 1214 VSS VSS nch l=0.26u w=0.8u
m2686 VSS 1217 VSS VSS nch l=0.26u w=0.8u
m2687 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2688 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2689 1297 1283 69923 VSS nch l=0.04u w=0.8u
m2690 69934 1290 VSS VSS nch l=0.04u w=0.8u
m2691 69935 1291 VSS VSS nch l=0.04u w=0.8u
m2692 VSS 1319 69924 VSS nch l=0.04u w=0.12u
m2693 VSS 1320 69925 VSS nch l=0.04u w=0.12u
m2694 1152 1353 1313 VSS nch l=0.04u w=0.4u
m2695 1312 1318 1280 VSS nch l=0.04u w=0.4u
m2696 69936 1438 1314 VSS nch l=0.04u w=0.8u
m2697 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2698 VSS 1229 VSS VSS nch l=0.26u w=0.8u
m2699 VSS 1230 VSS VSS nch l=0.26u w=0.8u
m2700 VSS 1233 VSS VSS nch l=0.26u w=0.8u
m2701 VSS 1235 VSS VSS nch l=0.26u w=0.8u
m2702 VSS 1236 VSS VSS nch l=0.26u w=0.8u
m2703 VSS 1239 VSS VSS nch l=0.26u w=0.8u
m2704 VSS 1372 1315 VSS nch l=0.04u w=0.4u
m2705 69937 977 69934 VSS nch l=0.04u w=0.8u
m2706 69938 978 69935 VSS nch l=0.04u w=0.8u
m2707 1319 1292 VSS VSS nch l=0.04u w=0.4u
m2708 1320 1293 VSS VSS nch l=0.04u w=0.4u
m2709 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2710 69939 1298 VSS VSS nch l=0.04u w=0.8u
m2711 1190 1336 272 VSS nch l=0.04u w=0.4u
m2712 69940 1299 VSS VSS nch l=0.04u w=0.8u
m2713 69941 1300 VSS VSS nch l=0.04u w=0.8u
m2714 1191 1337 139 VSS nch l=0.04u w=0.4u
m2715 69942 1301 VSS VSS nch l=0.04u w=0.8u
m2716 69943 1302 VSS VSS nch l=0.04u w=0.8u
m2717 1192 1338 FRAC[20] VSS nch l=0.04u w=0.4u
m2718 69944 1304 VSS VSS nch l=0.04u w=0.8u
m2719 1193 1341 960 VSS nch l=0.04u w=0.4u
m2720 69945 1305 VSS VSS nch l=0.04u w=0.8u
m2721 69946 1306 VSS VSS nch l=0.04u w=0.8u
m2722 1194 1342 820 VSS nch l=0.04u w=0.4u
m2723 69947 1307 VSS VSS nch l=0.04u w=0.8u
m2724 69948 1308 VSS VSS nch l=0.04u w=0.8u
m2725 69949 1309 VSS VSS nch l=0.04u w=0.8u
m2726 1195 1343 FRAC[20] VSS nch l=0.04u w=0.4u
m2727 69950 1310 VSS VSS nch l=0.04u w=0.8u
m2728 69951 1311 VSS VSS nch l=0.04u w=0.8u
m2729 VSS 1209 VSS VSS nch l=0.26u w=0.8u
m2730 VSS 1212 VSS VSS nch l=0.26u w=0.8u
m2731 VSS 1214 VSS VSS nch l=0.26u w=0.8u
m2732 VSS 1217 VSS VSS nch l=0.26u w=0.8u
m2733 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2734 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2735 1318 1280 1312 VSS nch l=0.04u w=0.4u
m2736 VSS 1394 69936 VSS nch l=0.04u w=0.8u
m2737 1335 1297 VSS VSS nch l=0.04u w=0.4u
m2738 1316 110 69937 VSS nch l=0.04u w=0.8u
m2739 1317 293 69938 VSS nch l=0.04u w=0.8u
m2740 69953 1003 69939 VSS nch l=0.04u w=0.8u
m2741 1336 272 1190 VSS nch l=0.04u w=0.4u
m2742 69954 1005 69940 VSS nch l=0.04u w=0.8u
m2743 69955 1006 69941 VSS nch l=0.04u w=0.8u
m2744 1337 139 1191 VSS nch l=0.04u w=0.4u
m2745 69956 1008 69942 VSS nch l=0.04u w=0.8u
m2746 69957 1009 69943 VSS nch l=0.04u w=0.8u
m2747 1338 FRAC[20] 1192 VSS nch l=0.04u w=0.4u
m2748 69958 1011 69944 VSS nch l=0.04u w=0.8u
m2749 1341 960 1193 VSS nch l=0.04u w=0.4u
m2750 69959 1014 69945 VSS nch l=0.04u w=0.8u
m2751 69960 1015 69946 VSS nch l=0.04u w=0.8u
m2752 1342 820 1194 VSS nch l=0.04u w=0.4u
m2753 69961 1017 69947 VSS nch l=0.04u w=0.8u
m2754 69962 1018 69948 VSS nch l=0.04u w=0.8u
m2755 69963 1019 69949 VSS nch l=0.04u w=0.8u
m2756 1343 FRAC[20] 1195 VSS nch l=0.04u w=0.4u
m2757 69964 1021 69950 VSS nch l=0.04u w=0.8u
m2758 69965 1022 69951 VSS nch l=0.04u w=0.8u
m2759 1346 1345 VSS VSS nch l=0.04u w=0.8u
m2760 1347 1348 VSS VSS nch l=0.04u w=0.8u
m2761 1350 1349 VSS VSS nch l=0.04u w=0.8u
m2762 1351 1352 VSS VSS nch l=0.04u w=0.8u
m2763 1353 1392 VSS VSS nch l=0.04u w=0.4u
m2764 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2765 VSS 1229 VSS VSS nch l=0.26u w=0.8u
m2766 VSS 1230 VSS VSS nch l=0.26u w=0.8u
m2767 VSS 1233 VSS VSS nch l=0.26u w=0.8u
m2768 VSS 1235 VSS VSS nch l=0.26u w=0.8u
m2769 VSS 1236 VSS VSS nch l=0.26u w=0.8u
m2770 VSS 1239 VSS VSS nch l=0.26u w=0.8u
m2771 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2772 VSS 1034 1296 VSS nch l=0.04u w=0.4u
m2773 1322 21 69953 VSS nch l=0.04u w=0.8u
m2774 VSS 1179 1336 VSS nch l=0.04u w=0.4u
m2775 1323 110 69954 VSS nch l=0.04u w=0.8u
m2776 1324 22 69955 VSS nch l=0.04u w=0.8u
m2777 VSS 1184 1337 VSS nch l=0.04u w=0.4u
m2778 1325 313 69956 VSS nch l=0.04u w=0.8u
m2779 1326 25 69957 VSS nch l=0.04u w=0.8u
m2780 VSS 94 1338 VSS nch l=0.04u w=0.4u
m2781 1327 315 69958 VSS nch l=0.04u w=0.8u
m2782 VSS 1319 1339 VSS nch l=0.04u w=0.4u
m2783 VSS 1320 1340 VSS nch l=0.04u w=0.4u
m2784 VSS 1321 1341 VSS nch l=0.04u w=0.4u
m2785 1328 27 69959 VSS nch l=0.04u w=0.8u
m2786 1329 28 69960 VSS nch l=0.04u w=0.8u
m2787 VSS 960 1342 VSS nch l=0.04u w=0.4u
m2788 1330 131 69961 VSS nch l=0.04u w=0.8u
m2789 1331 318 69962 VSS nch l=0.04u w=0.8u
m2790 1332 29 69963 VSS nch l=0.04u w=0.8u
m2791 VSS 961 1343 VSS nch l=0.04u w=0.4u
m2792 1333 131 69964 VSS nch l=0.04u w=0.8u
m2793 1334 318 69965 VSS nch l=0.04u w=0.8u
m2794 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2795 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2796 1356 377 VSS VSS nch l=0.04u w=0.4u
m2797 69967 REFDIV[5] 1354 VSS nch l=0.04u w=0.8u
m2798 1357 1358 VSS VSS nch l=0.04u w=0.8u
m2799 1360 1359 VSS VSS nch l=0.04u w=0.8u
m2800 1361 1362 VSS VSS nch l=0.04u w=0.8u
m2801 1363 1364 VSS VSS nch l=0.04u w=0.8u
m2802 1366 1365 VSS VSS nch l=0.04u w=0.8u
m2803 1367 1368 VSS VSS nch l=0.04u w=0.8u
m2804 69969 1511 VSS VSS nch l=0.04u w=0.8u
m2805 69970 1226 VSS VSS nch l=0.04u w=0.8u
m2806 69971 1227 VSS VSS nch l=0.04u w=0.8u
m2807 1001 1339 VSS VSS nch l=0.04u w=0.4u
m2808 793 1340 VSS VSS nch l=0.04u w=0.4u
m2809 VSS 1392 1355 VSS nch l=0.04u w=0.4u
m2810 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2811 VSS 377 69967 VSS nch l=0.04u w=0.8u
m2812 VSS 1178 VSS VSS nch l=0.26u w=0.8u
m2813 1369 1372 69969 VSS nch l=0.04u w=0.8u
m2814 1370 1316 69970 VSS nch l=0.04u w=0.8u
m2815 1371 1317 69971 VSS nch l=0.04u w=0.8u
m2816 VSS 1404 1372 VSS nch l=0.04u w=0.4u
m2817 69972 1242 VSS VSS nch l=0.04u w=0.8u
m2818 69973 1179 1373 VSS nch l=0.04u w=0.8u
m2819 69974 1243 VSS VSS nch l=0.04u w=0.8u
m2820 69975 1244 VSS VSS nch l=0.04u w=0.8u
m2821 69976 1184 1374 VSS nch l=0.04u w=0.8u
m2822 69977 1245 VSS VSS nch l=0.04u w=0.8u
m2823 69978 1246 VSS VSS nch l=0.04u w=0.8u
m2824 69979 94 1375 VSS nch l=0.04u w=0.8u
m2825 69980 1247 VSS VSS nch l=0.04u w=0.8u
m2826 69981 1321 1376 VSS nch l=0.04u w=0.8u
m2827 69982 1250 VSS VSS nch l=0.04u w=0.8u
m2828 69983 1251 VSS VSS nch l=0.04u w=0.8u
m2829 69984 960 1377 VSS nch l=0.04u w=0.8u
m2830 69985 1252 VSS VSS nch l=0.04u w=0.8u
m2831 69986 1253 VSS VSS nch l=0.04u w=0.8u
m2832 69987 1254 VSS VSS nch l=0.04u w=0.8u
m2833 69988 961 1378 VSS nch l=0.04u w=0.8u
m2834 69989 1255 VSS VSS nch l=0.04u w=0.8u
m2835 69990 1256 VSS VSS nch l=0.04u w=0.8u
m2836 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2837 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2838 69997 377 VSS VSS nch l=0.04u w=0.8u
m2839 1395 1396 VSS VSS nch l=0.04u w=0.8u
m2840 69998 1372 VSS VSS nch l=0.04u w=0.12u
m2841 1379 1322 69972 VSS nch l=0.04u w=0.8u
m2842 VSS 272 69973 VSS nch l=0.04u w=0.8u
m2843 1380 1323 69974 VSS nch l=0.04u w=0.8u
m2844 1381 1324 69975 VSS nch l=0.04u w=0.8u
m2845 VSS 139 69976 VSS nch l=0.04u w=0.8u
m2846 1382 1325 69977 VSS nch l=0.04u w=0.8u
m2847 1383 1326 69978 VSS nch l=0.04u w=0.8u
m2848 VSS FRAC[20] 69979 VSS nch l=0.04u w=0.8u
m2849 1384 1327 69980 VSS nch l=0.04u w=0.8u
m2850 1397 4328 VSS VSS nch l=0.04u w=0.4u
m2851 1398 4328 VSS VSS nch l=0.04u w=0.4u
m2852 VSS 960 69981 VSS nch l=0.04u w=0.8u
m2853 1385 1328 69982 VSS nch l=0.04u w=0.8u
m2854 1386 1329 69983 VSS nch l=0.04u w=0.8u
m2855 VSS 820 69984 VSS nch l=0.04u w=0.8u
m2856 1387 1330 69985 VSS nch l=0.04u w=0.8u
m2857 1388 1331 69986 VSS nch l=0.04u w=0.8u
m2858 1389 1332 69987 VSS nch l=0.04u w=0.8u
m2859 VSS FRAC[20] 69988 VSS nch l=0.04u w=0.8u
m2860 1390 1333 69989 VSS nch l=0.04u w=0.8u
m2861 1391 1334 69990 VSS nch l=0.04u w=0.8u
m2862 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2863 70003 1436 1392 VSS nch l=0.04u w=0.8u
m2864 1393 REFDIV[2] 69997 VSS nch l=0.04u w=0.8u
m2865 VSS 377 1394 VSS nch l=0.04u w=0.4u
m2866 1404 1529 69998 VSS nch l=0.04u w=0.12u
m2867 1401 1511 VSS VSS nch l=0.04u w=0.4u
m2868 VSS 1219 VSS VSS nch l=0.26u w=0.8u
m2869 VSS 1222 VSS VSS nch l=0.26u w=0.8u
m2870 70007 346 VSS VSS nch l=0.04u w=0.8u
m2871 70008 1447 VSS VSS nch l=0.04u w=0.8u
m2872 VSS 2648 70003 VSS nch l=0.04u w=0.8u
m2873 VSS 1399 1399 VSS nch l=0.04u w=0.8u
m2874 1412 1772 1404 VSS nch l=0.04u w=0.4u
m2875 VSS 1372 1401 VSS nch l=0.04u w=0.4u
m2876 1414 1413 VSS VSS nch l=0.04u w=0.8u
m2877 1415 1416 VSS VSS nch l=0.04u w=0.8u
m2878 1402 1179 70007 VSS nch l=0.04u w=0.8u
m2879 1403 129 70008 VSS nch l=0.04u w=0.8u
m2880 VSS 1405 1405 VSS nch l=0.04u w=0.8u
m2881 70010 1456 1159 VSS nch l=0.04u w=0.8u
m2882 70011 1503 VSS VSS nch l=0.04u w=0.8u
m2883 70012 1457 1162 VSS nch l=0.04u w=0.8u
m2884 70013 1514 VSS VSS nch l=0.04u w=0.8u
m2885 70014 2616 VSS VSS nch l=0.04u w=0.8u
m2886 70015 2616 VSS VSS nch l=0.04u w=0.8u
m2887 VSS 1407 1407 VSS nch l=0.04u w=0.8u
m2888 70016 2616 VSS VSS nch l=0.04u w=0.8u
m2889 70017 1458 1165 VSS nch l=0.04u w=0.8u
m2890 70018 FRAC[4] VSS VSS nch l=0.04u w=0.8u
m2891 1417 1397 1319 VSS nch l=0.04u w=0.4u
m2892 1418 1398 1320 VSS nch l=0.04u w=0.4u
m2893 VSS 1483 1409 VSS nch l=0.04u w=0.4u
m2894 70019 1504 VSS VSS nch l=0.04u w=0.8u
m2895 1426 4328 VSS VSS nch l=0.04u w=0.4u
m2896 1427 4328 VSS VSS nch l=0.04u w=0.4u
m2897 70020 1518 VSS VSS nch l=0.04u w=0.8u
m2898 70021 1460 1169 VSS nch l=0.04u w=0.8u
m2899 70022 1519 VSS VSS nch l=0.04u w=0.8u
m2900 70023 1409 VSS VSS nch l=0.04u w=0.8u
m2901 1431 4328 VSS VSS nch l=0.04u w=0.4u
m2902 1432 4328 VSS VSS nch l=0.04u w=0.4u
m2903 70024 1522 VSS VSS nch l=0.04u w=0.8u
m2904 70025 1461 1173 VSS nch l=0.04u w=0.8u
m2905 70026 FRAC[4] VSS VSS nch l=0.04u w=0.8u
m2906 70027 1409 VSS VSS nch l=0.04u w=0.8u
m2907 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2908 70028 1356 VSS VSS nch l=0.04u w=0.8u
m2909 1438 1448 1090 VSS nch l=0.04u w=0.4u
m2910 VSS 1411 1411 VSS nch l=0.04u w=0.8u
m2911 VSS 1618 70010 VSS nch l=0.04u w=0.8u
m2912 1419 1499 70011 VSS nch l=0.04u w=0.8u
m2913 VSS 1619 70012 VSS nch l=0.04u w=0.8u
m2914 1420 1502 70013 VSS nch l=0.04u w=0.8u
m2915 1421 1658 70014 VSS nch l=0.04u w=0.8u
m2916 1422 1659 70015 VSS nch l=0.04u w=0.8u
m2917 1423 1181 70016 VSS nch l=0.04u w=0.8u
m2918 VSS 1620 70017 VSS nch l=0.04u w=0.8u
m2919 1424 1503 70018 VSS nch l=0.04u w=0.8u
m2920 70030 4328 1417 VSS nch l=0.04u w=0.12u
m2921 70031 4328 1418 VSS nch l=0.04u w=0.12u
m2922 1425 131 70019 VSS nch l=0.04u w=0.8u
m2923 1428 1504 70020 VSS nch l=0.04u w=0.8u
m2924 VSS 1621 70021 VSS nch l=0.04u w=0.8u
m2925 1429 1505 70022 VSS nch l=0.04u w=0.8u
m2926 1430 1506 70023 VSS nch l=0.04u w=0.8u
m2927 1433 1507 70024 VSS nch l=0.04u w=0.8u
m2928 VSS 1622 70025 VSS nch l=0.04u w=0.8u
m2929 1434 1508 70026 VSS nch l=0.04u w=0.8u
m2930 1435 FBDIV[4] 70027 VSS nch l=0.04u w=0.8u
m2931 VSS 1484 1436 VSS nch l=0.04u w=0.4u
m2932 1437 1312 70028 VSS nch l=0.04u w=0.8u
m2933 1448 1090 1438 VSS nch l=0.04u w=0.4u
m2934 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m2935 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m2936 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m2937 VSS 1486 1412 VSS nch l=0.04u w=0.4u
m2938 1449 1335 VSS VSS nch l=0.04u w=0.4u
m2939 VSS 1440 1440 VSS nch l=0.04u w=0.8u
m2940 VSS 1441 1441 VSS nch l=0.04u w=0.8u
m2941 1450 1179 VSS VSS nch l=0.04u w=0.4u
m2942 1451 129 VSS VSS nch l=0.04u w=0.4u
m2943 VSS 1466 70030 VSS nch l=0.04u w=0.12u
m2944 VSS 1467 70031 VSS nch l=0.04u w=0.12u
m2945 1459 4328 VSS VSS nch l=0.04u w=0.4u
m2946 1452 1426 1443 VSS nch l=0.04u w=0.4u
m2947 1453 1427 1444 VSS nch l=0.04u w=0.4u
m2948 1454 1431 1445 VSS nch l=0.04u w=0.4u
m2949 1455 1432 1446 VSS nch l=0.04u w=0.4u
m2950 VSS 1264 VSS VSS nch l=0.26u w=0.8u
m2951 VSS 2906 1447 VSS nch l=0.04u w=0.4u
m2952 70035 1355 VSS VSS nch l=0.04u w=0.12u
m2953 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m2954 70036 1412 VSS VSS nch l=0.04u w=0.12u
m2955 1464 346 1450 VSS nch l=0.04u w=0.4u
m2956 1465 1447 1451 VSS nch l=0.04u w=0.4u
m2957 1466 1417 VSS VSS nch l=0.04u w=0.4u
m2958 1467 1418 VSS VSS nch l=0.04u w=0.4u
m2959 70037 2466 1456 VSS nch l=0.04u w=0.8u
m2960 1468 1499 VSS VSS nch l=0.04u w=0.4u
m2961 70038 2468 1457 VSS nch l=0.04u w=0.8u
m2962 1469 1502 VSS VSS nch l=0.04u w=0.4u
m2963 1470 1421 VSS VSS nch l=0.04u w=0.4u
m2964 1471 1422 VSS VSS nch l=0.04u w=0.4u
m2965 1472 1423 VSS VSS nch l=0.04u w=0.4u
m2966 70039 2470 1458 VSS nch l=0.04u w=0.8u
m2967 1473 1503 VSS VSS nch l=0.04u w=0.4u
m2968 1474 131 VSS VSS nch l=0.04u w=0.4u
m2969 70040 4328 1452 VSS nch l=0.04u w=0.12u
m2970 70041 4328 1453 VSS nch l=0.04u w=0.12u
m2971 1475 1504 VSS VSS nch l=0.04u w=0.4u
m2972 70042 2474 1460 VSS nch l=0.04u w=0.8u
m2973 1476 1505 VSS VSS nch l=0.04u w=0.4u
m2974 1477 1506 VSS VSS nch l=0.04u w=0.4u
m2975 70043 4328 1454 VSS nch l=0.04u w=0.12u
m2976 70044 4328 1455 VSS nch l=0.04u w=0.12u
m2977 1478 1507 VSS VSS nch l=0.04u w=0.4u
m2978 70045 2478 1461 VSS nch l=0.04u w=0.8u
m2979 1479 1508 VSS VSS nch l=0.04u w=0.4u
m2980 1480 FBDIV[4] VSS VSS nch l=0.04u w=0.4u
m2981 1482 1481 VSS VSS nch l=0.04u w=0.8u
m2982 1484 1623 70035 VSS nch l=0.04u w=0.12u
m2983 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m2984 70047 1437 VSS VSS nch l=0.04u w=0.8u
m2985 VSS 1448 1463 VSS nch l=0.04u w=0.4u
m2986 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m2987 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m2988 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m2989 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m2990 1486 1772 70036 VSS nch l=0.04u w=0.12u
m2991 346 1450 1464 VSS nch l=0.04u w=0.4u
m2992 1447 1451 1465 VSS nch l=0.04u w=0.4u
m2993 1487 1369 VSS VSS nch l=0.04u w=0.4u
m2994 70048 1671 70037 VSS nch l=0.04u w=0.8u
m2995 1488 1503 1468 VSS nch l=0.04u w=0.4u
m2996 70049 1672 70038 VSS nch l=0.04u w=0.8u
m2997 1489 1514 1469 VSS nch l=0.04u w=0.4u
m2998 70050 1673 70039 VSS nch l=0.04u w=0.8u
m2999 1490 FRAC[4] 1473 VSS nch l=0.04u w=0.4u
m3000 1492 1504 1474 VSS nch l=0.04u w=0.4u
m3001 VSS 1516 70040 VSS nch l=0.04u w=0.12u
m3002 VSS 1517 70041 VSS nch l=0.04u w=0.12u
m3003 1493 1518 1475 VSS nch l=0.04u w=0.4u
m3004 70051 1674 70042 VSS nch l=0.04u w=0.8u
m3005 1494 1519 1476 VSS nch l=0.04u w=0.4u
m3006 1495 1409 1477 VSS nch l=0.04u w=0.4u
m3007 VSS 1520 70043 VSS nch l=0.04u w=0.12u
m3008 VSS 1521 70044 VSS nch l=0.04u w=0.12u
m3009 1496 1522 1478 VSS nch l=0.04u w=0.4u
m3010 70052 1675 70045 VSS nch l=0.04u w=0.8u
m3011 1497 FRAC[4] 1479 VSS nch l=0.04u w=0.4u
m3012 1498 1409 1480 VSS nch l=0.04u w=0.4u
m3013 1491 1459 1483 VSS nch l=0.04u w=0.4u
m3014 1510 1663 1484 VSS nch l=0.04u w=0.4u
m3015 1485 1393 70047 VSS nch l=0.04u w=0.8u
m3016 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m3017 1511 1529 1486 VSS nch l=0.04u w=0.4u
m3018 VSS 1449 1487 VSS nch l=0.04u w=0.4u
m3019 VSS 1531 70048 VSS nch l=0.04u w=0.8u
m3020 1503 1468 1488 VSS nch l=0.04u w=0.4u
m3021 VSS 1533 70049 VSS nch l=0.04u w=0.8u
m3022 1514 1469 1489 VSS nch l=0.04u w=0.4u
m3023 VSS 1534 70050 VSS nch l=0.04u w=0.8u
m3024 FRAC[4] 1473 1490 VSS nch l=0.04u w=0.4u
m3025 1512 4328 1466 VSS nch l=0.04u w=0.4u
m3026 1513 4328 1467 VSS nch l=0.04u w=0.4u
m3027 1504 1474 1492 VSS nch l=0.04u w=0.4u
m3028 1516 1452 VSS VSS nch l=0.04u w=0.4u
m3029 1517 1453 VSS VSS nch l=0.04u w=0.4u
m3030 1518 1475 1493 VSS nch l=0.04u w=0.4u
m3031 VSS 1535 70051 VSS nch l=0.04u w=0.8u
m3032 1519 1476 1494 VSS nch l=0.04u w=0.4u
m3033 1409 1477 1495 VSS nch l=0.04u w=0.4u
m3034 1520 1454 VSS VSS nch l=0.04u w=0.4u
m3035 1521 1455 VSS VSS nch l=0.04u w=0.4u
m3036 1522 1478 1496 VSS nch l=0.04u w=0.4u
m3037 VSS 1536 70052 VSS nch l=0.04u w=0.8u
m3038 FRAC[4] 1479 1497 VSS nch l=0.04u w=0.4u
m3039 1409 1480 1498 VSS nch l=0.04u w=0.4u
m3040 1523 4328 VSS VSS nch l=0.04u w=0.4u
m3041 1524 4328 VSS VSS nch l=0.04u w=0.4u
m3042 1525 4328 VSS VSS nch l=0.04u w=0.4u
m3043 VSS 1501 1501 VSS nch l=0.04u w=0.8u
m3044 1526 4328 VSS VSS nch l=0.04u w=0.4u
m3045 1527 4328 VSS VSS nch l=0.04u w=0.4u
m3046 1528 4328 VSS VSS nch l=0.04u w=0.4u
m3047 70054 4328 1491 VSS nch l=0.04u w=0.12u
m3048 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m3049 70057 1393 1485 VSS nch l=0.04u w=0.8u
m3050 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m3051 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m3052 70058 683 1448 VSS nch l=0.04u w=0.8u
m3053 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m3054 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m3055 70059 1397 1512 VSS nch l=0.04u w=0.12u
m3056 70060 1398 1513 VSS nch l=0.04u w=0.12u
m3057 VSS 1550 70054 VSS nch l=0.04u w=0.12u
m3058 70072 1572 1510 VSS nch l=0.04u w=0.8u
m3059 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m3060 VSS 1437 70057 VSS nch l=0.04u w=0.8u
m3061 VSS 1561 70058 VSS nch l=0.04u w=0.8u
m3062 VSS 1772 1529 VSS nch l=0.04u w=0.4u
m3063 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3064 VSS 1562 70059 VSS nch l=0.04u w=0.12u
m3065 VSS 1563 70060 VSS nch l=0.04u w=0.12u
m3066 70073 1401 VSS VSS nch l=0.04u w=0.8u
m3067 70074 1464 1530 VSS nch l=0.04u w=0.8u
m3068 VSS 1564 1531 VSS nch l=0.04u w=0.4u
m3069 70075 1465 1532 VSS nch l=0.04u w=0.8u
m3070 VSS 1565 1533 VSS nch l=0.04u w=0.4u
m3071 VSS 1566 1534 VSS nch l=0.04u w=0.4u
m3072 1550 1491 VSS VSS nch l=0.04u w=0.4u
m3073 1539 4328 1516 VSS nch l=0.04u w=0.4u
m3074 1540 4328 1517 VSS nch l=0.04u w=0.4u
m3075 VSS 1567 1535 VSS nch l=0.04u w=0.4u
m3076 1541 4328 1520 VSS nch l=0.04u w=0.4u
m3077 1542 4328 1521 VSS nch l=0.04u w=0.4u
m3078 VSS 1568 1536 VSS nch l=0.04u w=0.4u
m3079 1544 1523 1537 VSS nch l=0.04u w=0.4u
m3080 1545 1524 1538 VSS nch l=0.04u w=0.4u
m3081 1546 1525 1180 VSS nch l=0.04u w=0.4u
m3082 1547 1526 1470 VSS nch l=0.04u w=0.4u
m3083 1548 1527 1471 VSS nch l=0.04u w=0.4u
m3084 1549 1528 1472 VSS nch l=0.04u w=0.4u
m3085 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m3086 VSS 2648 70072 VSS nch l=0.04u w=0.8u
m3087 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m3088 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m3089 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m3090 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m3091 1562 1512 VSS VSS nch l=0.04u w=0.4u
m3092 1563 1513 VSS VSS nch l=0.04u w=0.4u
m3093 1543 1335 70073 VSS nch l=0.04u w=0.8u
m3094 VSS 1370 70074 VSS nch l=0.04u w=0.8u
m3095 VSS 1371 70075 VSS nch l=0.04u w=0.8u
m3096 70076 1426 1539 VSS nch l=0.04u w=0.12u
m3097 70077 1427 1540 VSS nch l=0.04u w=0.12u
m3098 70078 1431 1541 VSS nch l=0.04u w=0.12u
m3099 70079 1432 1542 VSS nch l=0.04u w=0.12u
m3100 70080 4328 1544 VSS nch l=0.04u w=0.12u
m3101 70081 4328 1545 VSS nch l=0.04u w=0.12u
m3102 70082 4328 1546 VSS nch l=0.04u w=0.12u
m3103 70083 1488 1551 VSS nch l=0.04u w=0.8u
m3104 70084 1489 1552 VSS nch l=0.04u w=0.8u
m3105 70085 4328 1547 VSS nch l=0.04u w=0.12u
m3106 70086 4328 1548 VSS nch l=0.04u w=0.12u
m3107 70087 4328 1549 VSS nch l=0.04u w=0.12u
m3108 70088 1490 1553 VSS nch l=0.04u w=0.8u
m3109 70089 1492 1554 VSS nch l=0.04u w=0.8u
m3110 70090 1493 1555 VSS nch l=0.04u w=0.8u
m3111 70091 1494 1556 VSS nch l=0.04u w=0.8u
m3112 70092 1495 1557 VSS nch l=0.04u w=0.8u
m3113 70093 1496 1558 VSS nch l=0.04u w=0.8u
m3114 70094 1497 1559 VSS nch l=0.04u w=0.8u
m3115 70095 1498 1560 VSS nch l=0.04u w=0.8u
m3116 1569 155 VSS VSS nch l=0.04u w=0.4u
m3117 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m3118 70096 1510 VSS VSS nch l=0.04u w=0.24u
m3119 1570 76 VSS VSS nch l=0.04u w=0.4u
m3120 VSS 1573 1561 VSS nch l=0.04u w=0.4u
m3121 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3122 VSS 1592 1511 VSS nch l=0.04u w=0.4u
m3123 VSS 1576 70076 VSS nch l=0.04u w=0.12u
m3124 VSS 1577 70077 VSS nch l=0.04u w=0.12u
m3125 VSS 1578 70078 VSS nch l=0.04u w=0.12u
m3126 VSS 1579 70079 VSS nch l=0.04u w=0.12u
m3127 VSS 1582 70080 VSS nch l=0.04u w=0.12u
m3128 VSS 1583 70081 VSS nch l=0.04u w=0.12u
m3129 VSS 1584 70082 VSS nch l=0.04u w=0.12u
m3130 70097 1957 1564 VSS nch l=0.04u w=0.8u
m3131 VSS 1380 70083 VSS nch l=0.04u w=0.8u
m3132 70098 1958 1565 VSS nch l=0.04u w=0.8u
m3133 VSS 1382 70084 VSS nch l=0.04u w=0.8u
m3134 VSS 1586 70085 VSS nch l=0.04u w=0.12u
m3135 VSS 1587 70086 VSS nch l=0.04u w=0.12u
m3136 VSS 1588 70087 VSS nch l=0.04u w=0.12u
m3137 70099 1959 1566 VSS nch l=0.04u w=0.8u
m3138 VSS 1384 70088 VSS nch l=0.04u w=0.8u
m3139 1571 4328 1550 VSS nch l=0.04u w=0.4u
m3140 VSS 1385 70089 VSS nch l=0.04u w=0.8u
m3141 VSS 1386 70090 VSS nch l=0.04u w=0.8u
m3142 70100 1960 1567 VSS nch l=0.04u w=0.8u
m3143 VSS 1387 70091 VSS nch l=0.04u w=0.8u
m3144 VSS 1388 70092 VSS nch l=0.04u w=0.8u
m3145 VSS 1389 70093 VSS nch l=0.04u w=0.8u
m3146 70101 1961 1568 VSS nch l=0.04u w=0.8u
m3147 VSS 1390 70094 VSS nch l=0.04u w=0.8u
m3148 VSS 1391 70095 VSS nch l=0.04u w=0.8u
m3149 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m3150 1572 1663 70096 VSS nch l=0.04u w=0.24u
m3151 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m3152 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m3153 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m3154 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m3155 70102 1511 VSS VSS nch l=0.04u w=0.12u
m3156 1574 4328 VSS VSS nch l=0.04u w=0.4u
m3157 1575 4328 VSS VSS nch l=0.04u w=0.4u
m3158 1576 1539 VSS VSS nch l=0.04u w=0.4u
m3159 1577 1540 VSS VSS nch l=0.04u w=0.4u
m3160 1578 1541 VSS VSS nch l=0.04u w=0.4u
m3161 1579 1542 VSS VSS nch l=0.04u w=0.4u
m3162 1580 1543 VSS VSS nch l=0.04u w=0.4u
m3163 70103 1530 VSS VSS nch l=0.04u w=0.8u
m3164 1582 1544 VSS VSS nch l=0.04u w=0.4u
m3165 1583 1545 VSS VSS nch l=0.04u w=0.4u
m3166 1584 1546 VSS VSS nch l=0.04u w=0.4u
m3167 70104 2239 70097 VSS nch l=0.04u w=0.8u
m3168 70105 1532 VSS VSS nch l=0.04u w=0.8u
m3169 70106 2240 70098 VSS nch l=0.04u w=0.8u
m3170 1586 1547 VSS VSS nch l=0.04u w=0.4u
m3171 1587 1548 VSS VSS nch l=0.04u w=0.4u
m3172 1588 1549 VSS VSS nch l=0.04u w=0.4u
m3173 70107 2241 70099 VSS nch l=0.04u w=0.8u
m3174 70108 1459 1571 VSS nch l=0.04u w=0.12u
m3175 70109 2242 70100 VSS nch l=0.04u w=0.8u
m3176 70110 2243 70101 VSS nch l=0.04u w=0.8u
m3177 70111 155 VSS VSS nch l=0.04u w=0.8u
m3178 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m3179 1392 1623 1572 VSS nch l=0.04u w=0.4u
m3180 1591 1570 1485 VSS nch l=0.04u w=0.4u
m3181 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3182 70112 1240 1573 VSS nch l=0.04u w=0.8u
m3183 1592 1696 70102 VSS nch l=0.04u w=0.12u
m3184 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m3185 1581 1402 70103 VSS nch l=0.04u w=0.8u
m3186 VSS 2496 70104 VSS nch l=0.04u w=0.8u
m3187 1585 1403 70105 VSS nch l=0.04u w=0.8u
m3188 VSS 2497 70106 VSS nch l=0.04u w=0.8u
m3189 VSS 2498 70107 VSS nch l=0.04u w=0.8u
m3190 VSS 1613 70108 VSS nch l=0.04u w=0.12u
m3191 VSS 2499 70109 VSS nch l=0.04u w=0.8u
m3192 VSS 2500 70110 VSS nch l=0.04u w=0.8u
m3193 70113 1551 VSS VSS nch l=0.04u w=0.8u
m3194 70114 1552 VSS VSS nch l=0.04u w=0.8u
m3195 70115 1553 VSS VSS nch l=0.04u w=0.8u
m3196 70116 1554 VSS VSS nch l=0.04u w=0.8u
m3197 70117 1555 VSS VSS nch l=0.04u w=0.8u
m3198 70118 1556 VSS VSS nch l=0.04u w=0.8u
m3199 70119 1557 VSS VSS nch l=0.04u w=0.8u
m3200 70120 1558 VSS VSS nch l=0.04u w=0.8u
m3201 70121 1559 VSS VSS nch l=0.04u w=0.8u
m3202 70122 1560 VSS VSS nch l=0.04u w=0.8u
m3203 1589 FBDIV[4] 70111 VSS nch l=0.04u w=0.8u
m3204 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m3205 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m3206 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m3207 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m3208 70123 76 1591 VSS nch l=0.04u w=0.12u
m3209 70124 2194 70112 VSS nch l=0.04u w=0.8u
m3210 1604 1772 1592 VSS nch l=0.04u w=0.4u
m3211 1605 1574 1562 VSS nch l=0.04u w=0.4u
m3212 1606 1575 1563 VSS nch l=0.04u w=0.4u
m3213 1613 1571 VSS VSS nch l=0.04u w=0.4u
m3214 1614 4328 VSS VSS nch l=0.04u w=0.4u
m3215 1615 4328 VSS VSS nch l=0.04u w=0.4u
m3216 1616 4328 VSS VSS nch l=0.04u w=0.4u
m3217 1617 4328 VSS VSS nch l=0.04u w=0.4u
m3218 VSS 1637 1593 VSS nch l=0.04u w=0.4u
m3219 1607 4328 1582 VSS nch l=0.04u w=0.4u
m3220 1608 4328 1583 VSS nch l=0.04u w=0.4u
m3221 1609 4328 1584 VSS nch l=0.04u w=0.4u
m3222 1594 1419 70113 VSS nch l=0.04u w=0.8u
m3223 1595 1420 70114 VSS nch l=0.04u w=0.8u
m3224 1610 4328 1586 VSS nch l=0.04u w=0.4u
m3225 1611 4328 1587 VSS nch l=0.04u w=0.4u
m3226 1612 4328 1588 VSS nch l=0.04u w=0.4u
m3227 1596 1424 70115 VSS nch l=0.04u w=0.8u
m3228 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m3229 1597 1425 70116 VSS nch l=0.04u w=0.8u
m3230 1598 1428 70117 VSS nch l=0.04u w=0.8u
m3231 1599 1429 70118 VSS nch l=0.04u w=0.8u
m3232 1600 1430 70119 VSS nch l=0.04u w=0.8u
m3233 1601 1433 70120 VSS nch l=0.04u w=0.8u
m3234 1602 1434 70121 VSS nch l=0.04u w=0.8u
m3235 1603 1435 70122 VSS nch l=0.04u w=0.8u
m3236 1623 1663 VSS VSS nch l=0.04u w=0.4u
m3237 VSS 1631 70123 VSS nch l=0.04u w=0.12u
m3238 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3239 VSS 1653 70124 VSS nch l=0.04u w=0.8u
m3240 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m3241 70125 4328 1605 VSS nch l=0.04u w=0.12u
m3242 70126 4328 1606 VSS nch l=0.04u w=0.12u
m3243 70127 1593 VSS VSS nch l=0.04u w=0.12u
m3244 1624 1464 VSS VSS nch l=0.04u w=0.4u
m3245 70128 1523 1607 VSS nch l=0.04u w=0.12u
m3246 70129 1524 1608 VSS nch l=0.04u w=0.12u
m3247 70130 1525 1609 VSS nch l=0.04u w=0.12u
m3248 VSS 1719 1618 VSS nch l=0.04u w=0.4u
m3249 1625 1465 VSS VSS nch l=0.04u w=0.4u
m3250 VSS 1721 1619 VSS nch l=0.04u w=0.4u
m3251 70131 1526 1610 VSS nch l=0.04u w=0.12u
m3252 70132 1527 1611 VSS nch l=0.04u w=0.12u
m3253 70133 1528 1612 VSS nch l=0.04u w=0.12u
m3254 VSS 1726 1620 VSS nch l=0.04u w=0.4u
m3255 VSS 1730 1621 VSS nch l=0.04u w=0.4u
m3256 VSS 1734 1622 VSS nch l=0.04u w=0.4u
m3257 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m3258 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m3259 70135 1569 VSS VSS nch l=0.04u w=0.8u
m3260 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m3261 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m3262 1631 1591 VSS VSS nch l=0.04u w=0.4u
m3263 VSS 1666 1604 VSS nch l=0.04u w=0.4u
m3264 VSS 1654 70125 VSS nch l=0.04u w=0.12u
m3265 VSS 1655 70126 VSS nch l=0.04u w=0.12u
m3266 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m3267 1637 1744 70127 VSS nch l=0.04u w=0.12u
m3268 1636 1370 1624 VSS nch l=0.04u w=0.4u
m3269 VSS 979 70128 VSS nch l=0.04u w=0.12u
m3270 VSS 1499 70129 VSS nch l=0.04u w=0.12u
m3271 VSS 1023 70130 VSS nch l=0.04u w=0.12u
m3272 138 1371 1625 VSS nch l=0.04u w=0.4u
m3273 VSS 1657 70131 VSS nch l=0.04u w=0.12u
m3274 VSS 1503 70132 VSS nch l=0.04u w=0.12u
m3275 VSS 1027 70133 VSS nch l=0.04u w=0.12u
m3276 1632 1614 1626 VSS nch l=0.04u w=0.4u
m3277 1633 1615 1627 VSS nch l=0.04u w=0.4u
m3278 1634 1616 1628 VSS nch l=0.04u w=0.4u
m3279 1635 1617 1506 VSS nch l=0.04u w=0.4u
m3280 1639 1488 VSS VSS nch l=0.04u w=0.4u
m3281 1641 1489 VSS VSS nch l=0.04u w=0.4u
m3282 1643 1490 VSS VSS nch l=0.04u w=0.4u
m3283 1644 1492 VSS VSS nch l=0.04u w=0.4u
m3284 1645 1493 VSS VSS nch l=0.04u w=0.4u
m3285 1647 1494 VSS VSS nch l=0.04u w=0.4u
m3286 1648 1495 VSS VSS nch l=0.04u w=0.4u
m3287 1649 1496 VSS VSS nch l=0.04u w=0.4u
m3288 1651 1497 VSS VSS nch l=0.04u w=0.4u
m3289 1652 1498 VSS VSS nch l=0.04u w=0.4u
m3290 1629 1613 70135 VSS nch l=0.04u w=0.8u
m3291 VSS 1663 1630 VSS nch l=0.04u w=0.4u
m3292 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3293 1653 1677 VSS VSS nch l=0.04u w=0.4u
m3294 VSS 1400 VSS VSS nch l=0.26u w=0.8u
m3295 70142 1604 VSS VSS nch l=0.04u w=0.12u
m3296 1654 1605 VSS VSS nch l=0.04u w=0.4u
m3297 1655 1606 VSS VSS nch l=0.04u w=0.4u
m3298 1656 3012 1637 VSS nch l=0.04u w=0.4u
m3299 1370 1624 1636 VSS nch l=0.04u w=0.4u
m3300 979 1607 VSS VSS nch l=0.04u w=0.4u
m3301 1499 1608 VSS VSS nch l=0.04u w=0.4u
m3302 VSS 1406 VSS VSS nch l=0.26u w=0.8u
m3303 1023 1609 VSS VSS nch l=0.04u w=0.4u
m3304 1371 1625 138 VSS nch l=0.04u w=0.4u
m3305 1657 1610 VSS VSS nch l=0.04u w=0.4u
m3306 1503 1611 VSS VSS nch l=0.04u w=0.4u
m3307 VSS 1408 VSS VSS nch l=0.26u w=0.8u
m3308 1027 1612 VSS VSS nch l=0.04u w=0.4u
m3309 70144 4328 1632 VSS nch l=0.04u w=0.12u
m3310 70145 4328 1633 VSS nch l=0.04u w=0.12u
m3311 70146 4328 1634 VSS nch l=0.04u w=0.12u
m3312 70147 4328 1635 VSS nch l=0.04u w=0.12u
m3313 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m3314 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m3315 1538 1380 1639 VSS nch l=0.04u w=0.4u
m3316 1659 1382 1641 VSS nch l=0.04u w=0.4u
m3317 1502 1384 1643 VSS nch l=0.04u w=0.4u
m3318 1483 1385 1644 VSS nch l=0.04u w=0.4u
m3319 1627 1386 1645 VSS nch l=0.04u w=0.4u
m3320 1661 1387 1647 VSS nch l=0.04u w=0.4u
m3321 1518 1388 1648 VSS nch l=0.04u w=0.4u
m3322 1506 1389 1649 VSS nch l=0.04u w=0.4u
m3323 1519 1390 1651 VSS nch l=0.04u w=0.4u
m3324 1522 1391 1652 VSS nch l=0.04u w=0.4u
m3325 1662 76 1631 VSS nch l=0.04u w=0.4u
m3326 VSS 1677 1653 VSS nch l=0.04u w=0.4u
m3327 1664 1665 VSS VSS nch l=0.04u w=0.8u
m3328 VSS 1410 VSS VSS nch l=0.26u w=0.8u
m3329 1666 1772 70142 VSS nch l=0.04u w=0.12u
m3330 1667 1668 VSS VSS nch l=0.04u w=0.8u
m3331 1669 1670 VSS VSS nch l=0.04u w=0.8u
m3332 VSS 1685 70144 VSS nch l=0.04u w=0.12u
m3333 VSS 1686 70145 VSS nch l=0.04u w=0.12u
m3334 VSS 1687 70146 VSS nch l=0.04u w=0.12u
m3335 VSS 1688 70147 VSS nch l=0.04u w=0.12u
m3336 1380 1639 1538 VSS nch l=0.04u w=0.4u
m3337 1382 1641 1659 VSS nch l=0.04u w=0.4u
m3338 1384 1643 1502 VSS nch l=0.04u w=0.4u
m3339 1385 1644 1483 VSS nch l=0.04u w=0.4u
m3340 1386 1645 1627 VSS nch l=0.04u w=0.4u
m3341 1387 1647 1661 VSS nch l=0.04u w=0.4u
m3342 1388 1648 1518 VSS nch l=0.04u w=0.4u
m3343 1389 1649 1506 VSS nch l=0.04u w=0.4u
m3344 1390 1651 1519 VSS nch l=0.04u w=0.4u
m3345 1391 1652 1522 VSS nch l=0.04u w=0.4u
m3346 1537 1689 1638 VSS nch l=0.04u w=0.4u
m3347 1658 1690 1640 VSS nch l=0.04u w=0.4u
m3348 1660 1691 1642 VSS nch l=0.04u w=0.4u
m3349 1444 1692 1646 VSS nch l=0.04u w=0.4u
m3350 1446 1693 1650 VSS nch l=0.04u w=0.4u
m3351 70149 1629 VSS VSS nch l=0.04u w=0.8u
m3352 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3353 70158 1708 1663 VSS nch l=0.04u w=0.8u
m3354 70159 1570 1662 VSS nch l=0.04u w=0.12u
m3355 1681 1680 VSS VSS nch l=0.04u w=0.8u
m3356 1682 1696 1666 VSS nch l=0.04u w=0.4u
m3357 VSS 1439 VSS VSS nch l=0.26u w=0.8u
m3358 VSS 1442 VSS VSS nch l=0.26u w=0.8u
m3359 1683 4328 1654 VSS nch l=0.04u w=0.4u
m3360 1684 4328 1655 VSS nch l=0.04u w=0.4u
m3361 1685 1632 VSS VSS nch l=0.04u w=0.4u
m3362 1686 1633 VSS VSS nch l=0.04u w=0.4u
m3363 1687 1634 VSS VSS nch l=0.04u w=0.4u
m3364 1688 1635 VSS VSS nch l=0.04u w=0.4u
m3365 VSS 1718 1656 VSS nch l=0.04u w=0.4u
m3366 1689 1638 1537 VSS nch l=0.04u w=0.4u
m3367 1690 1640 1658 VSS nch l=0.04u w=0.4u
m3368 1691 1642 1660 VSS nch l=0.04u w=0.4u
m3369 1692 1646 1444 VSS nch l=0.04u w=0.4u
m3370 1693 1650 1446 VSS nch l=0.04u w=0.4u
m3371 1676 1589 70149 VSS nch l=0.04u w=0.8u
m3372 VSS 2648 70158 VSS nch l=0.04u w=0.8u
m3373 VSS 1318 70159 VSS nch l=0.04u w=0.12u
m3374 VSS 1737 1677 VSS nch l=0.04u w=0.4u
m3375 VSS 1678 1678 VSS nch l=0.04u w=0.8u
m3376 1698 1697 VSS VSS nch l=0.04u w=0.8u
m3377 1699 1700 VSS VSS nch l=0.04u w=0.8u
m3378 70176 1574 1683 VSS nch l=0.04u w=0.12u
m3379 70177 1575 1684 VSS nch l=0.04u w=0.12u
m3380 70178 1656 VSS VSS nch l=0.04u w=0.12u
m3381 70182 110 VSS VSS nch l=0.04u w=0.8u
m3382 VSS 1671 1689 VSS nch l=0.04u w=0.4u
m3383 70183 1741 VSS VSS nch l=0.04u w=0.8u
m3384 VSS 1672 1690 VSS nch l=0.04u w=0.4u
m3385 VSS 1673 1691 VSS nch l=0.04u w=0.4u
m3386 VSS 1674 1692 VSS nch l=0.04u w=0.4u
m3387 VSS 1675 1693 VSS nch l=0.04u w=0.4u
m3388 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3389 1318 1662 VSS VSS nch l=0.04u w=0.4u
m3390 70184 1677 VSS VSS nch l=0.04u w=0.12u
m3391 VSS 1695 1695 VSS nch l=0.04u w=0.8u
m3392 VSS 1772 1696 VSS nch l=0.04u w=0.4u
m3393 VSS 1738 70176 VSS nch l=0.04u w=0.12u
m3394 VSS 1739 70177 VSS nch l=0.04u w=0.12u
m3395 1718 3012 70178 VSS nch l=0.04u w=0.12u
m3396 1710 4328 1685 VSS nch l=0.04u w=0.4u
m3397 1711 4328 1686 VSS nch l=0.04u w=0.4u
m3398 1712 4328 1687 VSS nch l=0.04u w=0.4u
m3399 1713 4328 1688 VSS nch l=0.04u w=0.4u
m3400 1701 888 70182 VSS nch l=0.04u w=0.8u
m3401 1702 441 70183 VSS nch l=0.04u w=0.8u
m3402 VSS 1703 1703 VSS nch l=0.04u w=0.8u
m3403 70187 1791 VSS VSS nch l=0.04u w=0.8u
m3404 70188 1803 VSS VSS nch l=0.04u w=0.8u
m3405 70189 2616 VSS VSS nch l=0.04u w=0.8u
m3406 70190 2616 VSS VSS nch l=0.04u w=0.8u
m3407 VSS 1705 1705 VSS nch l=0.04u w=0.8u
m3408 70191 2616 VSS VSS nch l=0.04u w=0.8u
m3409 70192 FRAC[5] VSS VSS nch l=0.04u w=0.8u
m3410 VSS 1770 1707 VSS nch l=0.04u w=0.4u
m3411 70193 1792 VSS VSS nch l=0.04u w=0.8u
m3412 70194 1805 VSS VSS nch l=0.04u w=0.8u
m3413 70195 1628 VSS VSS nch l=0.04u w=0.8u
m3414 70196 1707 VSS VSS nch l=0.04u w=0.8u
m3415 70197 1806 VSS VSS nch l=0.04u w=0.8u
m3416 70198 FRAC[5] VSS VSS nch l=0.04u w=0.8u
m3417 70199 1707 VSS VSS nch l=0.04u w=0.8u
m3418 VSS 1750 1708 VSS nch l=0.04u w=0.4u
m3419 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3420 1737 1844 70184 VSS nch l=0.04u w=0.12u
m3421 1738 1683 VSS VSS nch l=0.04u w=0.4u
m3422 1739 1684 VSS VSS nch l=0.04u w=0.4u
m3423 1740 1744 1718 VSS nch l=0.04u w=0.4u
m3424 VSS 1715 1715 VSS nch l=0.04u w=0.8u
m3425 VSS 1716 1716 VSS nch l=0.04u w=0.8u
m3426 70201 1614 1710 VSS nch l=0.04u w=0.12u
m3427 70202 1615 1711 VSS nch l=0.04u w=0.12u
m3428 70203 1616 1712 VSS nch l=0.04u w=0.12u
m3429 70204 1617 1713 VSS nch l=0.04u w=0.12u
m3430 VSS 1500 VSS VSS nch l=0.26u w=0.8u
m3431 70205 1879 1719 VSS nch l=0.04u w=0.8u
m3432 1720 1789 70187 VSS nch l=0.04u w=0.8u
m3433 70206 1881 1721 VSS nch l=0.04u w=0.8u
m3434 1722 1790 70188 VSS nch l=0.04u w=0.8u
m3435 1723 1944 70189 VSS nch l=0.04u w=0.8u
m3436 1724 1945 70190 VSS nch l=0.04u w=0.8u
m3437 1725 892 70191 VSS nch l=0.04u w=0.8u
m3438 70207 1883 1726 VSS nch l=0.04u w=0.8u
m3439 1727 1791 70192 VSS nch l=0.04u w=0.8u
m3440 1728 131 70193 VSS nch l=0.04u w=0.8u
m3441 1729 1792 70194 VSS nch l=0.04u w=0.8u
m3442 70208 1887 1730 VSS nch l=0.04u w=0.8u
m3443 1731 1753 70195 VSS nch l=0.04u w=0.8u
m3444 1732 1793 70196 VSS nch l=0.04u w=0.8u
m3445 1733 1794 70197 VSS nch l=0.04u w=0.8u
m3446 70209 1891 1734 VSS nch l=0.04u w=0.8u
m3447 1735 1754 70198 VSS nch l=0.04u w=0.8u
m3448 1736 FBDIV[5] 70199 VSS nch l=0.04u w=0.8u
m3449 70211 1630 VSS VSS nch l=0.04u w=0.12u
m3450 1742 1318 VSS VSS nch l=0.04u w=0.4u
m3451 1743 76 1737 VSS nch l=0.04u w=0.4u
m3452 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3453 VSS 1372 1682 VSS nch l=0.04u w=0.4u
m3454 VSS 1753 70201 VSS nch l=0.04u w=0.12u
m3455 VSS 1504 70202 VSS nch l=0.04u w=0.12u
m3456 VSS 1754 70203 VSS nch l=0.04u w=0.12u
m3457 VSS 1507 70204 VSS nch l=0.04u w=0.12u
m3458 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3459 1746 1745 VSS VSS nch l=0.04u w=0.8u
m3460 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3461 1747 888 VSS VSS nch l=0.04u w=0.4u
m3462 VSS 1773 70205 VSS nch l=0.04u w=0.8u
m3463 1748 441 VSS VSS nch l=0.04u w=0.4u
m3464 VSS 1775 70206 VSS nch l=0.04u w=0.8u
m3465 VSS 1777 70207 VSS nch l=0.04u w=0.8u
m3466 VSS 1782 70208 VSS nch l=0.04u w=0.8u
m3467 VSS 1786 70209 VSS nch l=0.04u w=0.8u
m3468 1749 4328 VSS VSS nch l=0.04u w=0.4u
m3469 VSS 3180 1741 VSS nch l=0.04u w=0.4u
m3470 1750 1894 70211 VSS nch l=0.04u w=0.12u
m3471 VSS 1318 1742 VSS nch l=0.04u w=0.4u
m3472 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3473 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3474 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3475 1751 4328 VSS VSS nch l=0.04u w=0.4u
m3476 1752 4328 VSS VSS nch l=0.04u w=0.4u
m3477 1753 1710 VSS VSS nch l=0.04u w=0.4u
m3478 1504 1711 VSS VSS nch l=0.04u w=0.4u
m3479 1754 1712 VSS VSS nch l=0.04u w=0.4u
m3480 1507 1713 VSS VSS nch l=0.04u w=0.4u
m3481 VSS 3012 1744 VSS nch l=0.04u w=0.4u
m3482 1755 110 1747 VSS nch l=0.04u w=0.4u
m3483 1756 1741 1748 VSS nch l=0.04u w=0.4u
m3484 1757 1789 VSS VSS nch l=0.04u w=0.4u
m3485 1758 1790 VSS VSS nch l=0.04u w=0.4u
m3486 1759 1723 VSS VSS nch l=0.04u w=0.4u
m3487 1760 1724 VSS VSS nch l=0.04u w=0.4u
m3488 1761 1725 VSS VSS nch l=0.04u w=0.4u
m3489 1762 1791 VSS VSS nch l=0.04u w=0.4u
m3490 1763 131 VSS VSS nch l=0.04u w=0.4u
m3491 1764 1792 VSS VSS nch l=0.04u w=0.4u
m3492 1765 1753 VSS VSS nch l=0.04u w=0.4u
m3493 1766 1793 VSS VSS nch l=0.04u w=0.4u
m3494 1767 1794 VSS VSS nch l=0.04u w=0.4u
m3495 1768 1754 VSS VSS nch l=0.04u w=0.4u
m3496 1769 FBDIV[5] VSS VSS nch l=0.04u w=0.4u
m3497 1771 1934 1750 VSS nch l=0.04u w=0.4u
m3498 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3499 VSS 1813 1743 VSS nch l=0.04u w=0.4u
m3500 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3501 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3502 1772 1848 VSS VSS nch l=0.04u w=0.4u
m3503 110 1747 1755 VSS nch l=0.04u w=0.4u
m3504 1741 1748 1756 VSS nch l=0.04u w=0.4u
m3505 70216 1638 VSS VSS nch l=0.04u w=0.8u
m3506 1774 1791 1757 VSS nch l=0.04u w=0.4u
m3507 70217 1640 VSS VSS nch l=0.04u w=0.8u
m3508 1776 1803 1758 VSS nch l=0.04u w=0.4u
m3509 70218 1642 VSS VSS nch l=0.04u w=0.8u
m3510 1778 FRAC[5] 1762 VSS nch l=0.04u w=0.4u
m3511 1780 1792 1763 VSS nch l=0.04u w=0.4u
m3512 1781 1805 1764 VSS nch l=0.04u w=0.4u
m3513 70219 1646 VSS VSS nch l=0.04u w=0.8u
m3514 1783 1628 1765 VSS nch l=0.04u w=0.4u
m3515 1784 1707 1766 VSS nch l=0.04u w=0.4u
m3516 1785 1806 1767 VSS nch l=0.04u w=0.4u
m3517 70220 1650 VSS VSS nch l=0.04u w=0.8u
m3518 1787 FRAC[5] 1768 VSS nch l=0.04u w=0.4u
m3519 1788 1707 1769 VSS nch l=0.04u w=0.4u
m3520 1779 1749 1770 VSS nch l=0.04u w=0.4u
m3521 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3522 70222 1742 VSS VSS nch l=0.04u w=0.8u
m3523 70223 1743 VSS VSS nch l=0.04u w=0.12u
m3524 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3525 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3526 VSS 1848 1772 VSS nch l=0.04u w=0.4u
m3527 1797 1751 1738 VSS nch l=0.04u w=0.4u
m3528 1798 1752 1739 VSS nch l=0.04u w=0.4u
m3529 1799 4328 VSS VSS nch l=0.04u w=0.4u
m3530 1800 4328 VSS VSS nch l=0.04u w=0.4u
m3531 1801 4328 VSS VSS nch l=0.04u w=0.4u
m3532 1802 4328 VSS VSS nch l=0.04u w=0.4u
m3533 VSS 1826 1740 VSS nch l=0.04u w=0.4u
m3534 1773 1671 70216 VSS nch l=0.04u w=0.8u
m3535 1791 1757 1774 VSS nch l=0.04u w=0.4u
m3536 1775 1672 70217 VSS nch l=0.04u w=0.8u
m3537 1803 1758 1776 VSS nch l=0.04u w=0.4u
m3538 1777 1673 70218 VSS nch l=0.04u w=0.8u
m3539 FRAC[5] 1762 1778 VSS nch l=0.04u w=0.4u
m3540 1792 1763 1780 VSS nch l=0.04u w=0.4u
m3541 1805 1764 1781 VSS nch l=0.04u w=0.4u
m3542 1782 1674 70219 VSS nch l=0.04u w=0.8u
m3543 1628 1765 1783 VSS nch l=0.04u w=0.4u
m3544 1707 1766 1784 VSS nch l=0.04u w=0.4u
m3545 1806 1767 1785 VSS nch l=0.04u w=0.4u
m3546 1786 1675 70220 VSS nch l=0.04u w=0.8u
m3547 FRAC[5] 1768 1787 VSS nch l=0.04u w=0.4u
m3548 1707 1769 1788 VSS nch l=0.04u w=0.4u
m3549 1807 4328 VSS VSS nch l=0.04u w=0.4u
m3550 1808 4328 VSS VSS nch l=0.04u w=0.4u
m3551 1809 4328 VSS VSS nch l=0.04u w=0.4u
m3552 1810 4328 VSS VSS nch l=0.04u w=0.4u
m3553 1811 4328 VSS VSS nch l=0.04u w=0.4u
m3554 1812 4328 VSS VSS nch l=0.04u w=0.4u
m3555 70224 4328 1779 VSS nch l=0.04u w=0.12u
m3556 70228 1851 1771 VSS nch l=0.04u w=0.8u
m3557 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3558 70229 1240 70222 VSS nch l=0.04u w=0.8u
m3559 1813 76 70223 VSS nch l=0.04u w=0.12u
m3560 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3561 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3562 1772 1848 VSS VSS nch l=0.04u w=0.4u
m3563 70231 4328 1797 VSS nch l=0.04u w=0.12u
m3564 70232 4328 1798 VSS nch l=0.04u w=0.12u
m3565 70234 1740 VSS VSS nch l=0.04u w=0.12u
m3566 VSS 1833 70224 VSS nch l=0.04u w=0.12u
m3567 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3568 VSS 2648 70228 VSS nch l=0.04u w=0.8u
m3569 1796 683 70229 VSS nch l=0.04u w=0.8u
m3570 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3571 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3572 1821 1844 1813 VSS nch l=0.04u w=0.4u
m3573 VSS 1848 1772 VSS nch l=0.04u w=0.4u
m3574 VSS 1846 70231 VSS nch l=0.04u w=0.12u
m3575 VSS 1847 70232 VSS nch l=0.04u w=0.12u
m3576 1826 1917 70234 VSS nch l=0.04u w=0.12u
m3577 1822 1799 1814 VSS nch l=0.04u w=0.4u
m3578 1823 1800 1661 VSS nch l=0.04u w=0.4u
m3579 1824 1801 1815 VSS nch l=0.04u w=0.4u
m3580 1825 1802 1519 VSS nch l=0.04u w=0.4u
m3581 70250 1755 1816 VSS nch l=0.04u w=0.8u
m3582 70251 1756 1817 VSS nch l=0.04u w=0.8u
m3583 1833 1779 VSS VSS nch l=0.04u w=0.4u
m3584 1827 1807 1819 VSS nch l=0.04u w=0.4u
m3585 1828 1808 1820 VSS nch l=0.04u w=0.4u
m3586 1829 1809 891 VSS nch l=0.04u w=0.4u
m3587 1830 1810 1759 VSS nch l=0.04u w=0.4u
m3588 1831 1811 1760 VSS nch l=0.04u w=0.4u
m3589 1832 1812 1761 VSS nch l=0.04u w=0.4u
m3590 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3591 70253 1771 VSS VSS nch l=0.04u w=0.24u
m3592 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3593 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3594 1846 1797 VSS VSS nch l=0.04u w=0.4u
m3595 1847 1798 VSS VSS nch l=0.04u w=0.4u
m3596 1849 3012 1826 VSS nch l=0.04u w=0.4u
m3597 70254 4328 1822 VSS nch l=0.04u w=0.12u
m3598 70255 4328 1823 VSS nch l=0.04u w=0.12u
m3599 70256 4328 1824 VSS nch l=0.04u w=0.12u
m3600 70257 4328 1825 VSS nch l=0.04u w=0.12u
m3601 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3602 VSS 1581 70250 VSS nch l=0.04u w=0.8u
m3603 VSS 1585 70251 VSS nch l=0.04u w=0.8u
m3604 70258 4328 1827 VSS nch l=0.04u w=0.12u
m3605 70259 4328 1828 VSS nch l=0.04u w=0.12u
m3606 70260 4328 1829 VSS nch l=0.04u w=0.12u
m3607 1671 1855 1657 VSS nch l=0.04u w=0.4u
m3608 70261 1774 1834 VSS nch l=0.04u w=0.8u
m3609 1672 1856 139 VSS nch l=0.04u w=0.4u
m3610 70262 1776 1835 VSS nch l=0.04u w=0.8u
m3611 70263 4328 1830 VSS nch l=0.04u w=0.12u
m3612 70264 4328 1831 VSS nch l=0.04u w=0.12u
m3613 70265 4328 1832 VSS nch l=0.04u w=0.12u
m3614 1673 1857 FRAC[19] VSS nch l=0.04u w=0.4u
m3615 70266 1778 1836 VSS nch l=0.04u w=0.8u
m3616 70267 1780 1837 VSS nch l=0.04u w=0.8u
m3617 70268 1781 1838 VSS nch l=0.04u w=0.8u
m3618 1674 1858 1446 VSS nch l=0.04u w=0.4u
m3619 70269 1783 1839 VSS nch l=0.04u w=0.8u
m3620 70270 1784 1840 VSS nch l=0.04u w=0.8u
m3621 70271 1785 1841 VSS nch l=0.04u w=0.8u
m3622 1675 1859 FRAC[19] VSS nch l=0.04u w=0.4u
m3623 70272 1787 1842 VSS nch l=0.04u w=0.8u
m3624 70273 1788 1843 VSS nch l=0.04u w=0.8u
m3625 1850 155 VSS VSS nch l=0.04u w=0.4u
m3626 1851 1934 70253 VSS nch l=0.04u w=0.24u
m3627 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3628 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3629 1852 1796 VSS VSS nch l=0.04u w=0.4u
m3630 1853 1943 VSS VSS nch l=0.04u w=0.4u
m3631 VSS 76 1844 VSS nch l=0.04u w=0.4u
m3632 70274 1916 1848 VSS nch l=0.04u w=0.8u
m3633 VSS 1863 70254 VSS nch l=0.04u w=0.12u
m3634 VSS 1864 70255 VSS nch l=0.04u w=0.12u
m3635 VSS 1865 70256 VSS nch l=0.04u w=0.12u
m3636 VSS 1866 70257 VSS nch l=0.04u w=0.12u
m3637 VSS 1868 70258 VSS nch l=0.04u w=0.12u
m3638 VSS 1869 70259 VSS nch l=0.04u w=0.12u
m3639 VSS 1870 70260 VSS nch l=0.04u w=0.12u
m3640 1855 1657 1671 VSS nch l=0.04u w=0.4u
m3641 VSS 1594 70261 VSS nch l=0.04u w=0.8u
m3642 1856 139 1672 VSS nch l=0.04u w=0.4u
m3643 VSS 1595 70262 VSS nch l=0.04u w=0.8u
m3644 VSS 1872 70263 VSS nch l=0.04u w=0.12u
m3645 VSS 1873 70264 VSS nch l=0.04u w=0.12u
m3646 VSS 1874 70265 VSS nch l=0.04u w=0.12u
m3647 1857 FRAC[19] 1673 VSS nch l=0.04u w=0.4u
m3648 VSS 1596 70266 VSS nch l=0.04u w=0.8u
m3649 1854 4328 1833 VSS nch l=0.04u w=0.4u
m3650 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3651 VSS 1597 70267 VSS nch l=0.04u w=0.8u
m3652 VSS 1598 70268 VSS nch l=0.04u w=0.8u
m3653 1858 1446 1674 VSS nch l=0.04u w=0.4u
m3654 VSS 1599 70269 VSS nch l=0.04u w=0.8u
m3655 VSS 1600 70270 VSS nch l=0.04u w=0.8u
m3656 VSS 1601 70271 VSS nch l=0.04u w=0.8u
m3657 1859 FRAC[19] 1675 VSS nch l=0.04u w=0.4u
m3658 VSS 1602 70272 VSS nch l=0.04u w=0.8u
m3659 VSS 1603 70273 VSS nch l=0.04u w=0.8u
m3660 1663 1894 1851 VSS nch l=0.04u w=0.4u
m3661 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3662 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3663 VSS 1878 70274 VSS nch l=0.04u w=0.8u
m3664 1861 4328 1846 VSS nch l=0.04u w=0.4u
m3665 1862 4328 1847 VSS nch l=0.04u w=0.4u
m3666 1863 1822 VSS VSS nch l=0.04u w=0.4u
m3667 1864 1823 VSS VSS nch l=0.04u w=0.4u
m3668 1865 1824 VSS VSS nch l=0.04u w=0.4u
m3669 1866 1825 VSS VSS nch l=0.04u w=0.4u
m3670 VSS 1899 1849 VSS nch l=0.04u w=0.4u
m3671 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3672 70275 1816 VSS VSS nch l=0.04u w=0.8u
m3673 1868 1827 VSS VSS nch l=0.04u w=0.4u
m3674 1869 1828 VSS VSS nch l=0.04u w=0.4u
m3675 1870 1829 VSS VSS nch l=0.04u w=0.4u
m3676 VSS 979 1855 VSS nch l=0.04u w=0.4u
m3677 70276 1817 VSS VSS nch l=0.04u w=0.8u
m3678 VSS 1660 1856 VSS nch l=0.04u w=0.4u
m3679 1872 1830 VSS VSS nch l=0.04u w=0.4u
m3680 1873 1831 VSS VSS nch l=0.04u w=0.4u
m3681 1874 1832 VSS VSS nch l=0.04u w=0.4u
m3682 VSS 1657 1857 VSS nch l=0.04u w=0.4u
m3683 70277 1749 1854 VSS nch l=0.04u w=0.12u
m3684 VSS 1577 1858 VSS nch l=0.04u w=0.4u
m3685 VSS 1579 1859 VSS nch l=0.04u w=0.4u
m3686 70278 155 VSS VSS nch l=0.04u w=0.8u
m3687 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3688 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3689 1860 1876 1796 VSS nch l=0.04u w=0.4u
m3690 1877 1657 VSS VSS nch l=0.04u w=0.4u
m3691 70279 1936 VSS VSS nch l=0.04u w=0.8u
m3692 70280 1751 1861 VSS nch l=0.04u w=0.12u
m3693 70281 1752 1862 VSS nch l=0.04u w=0.12u
m3694 70282 1849 VSS VSS nch l=0.04u w=0.12u
m3695 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3696 1867 1701 70275 VSS nch l=0.04u w=0.8u
m3697 1871 1702 70276 VSS nch l=0.04u w=0.8u
m3698 VSS 1906 70277 VSS nch l=0.04u w=0.12u
m3699 70283 1834 VSS VSS nch l=0.04u w=0.8u
m3700 70284 1835 VSS VSS nch l=0.04u w=0.8u
m3701 70285 1836 VSS VSS nch l=0.04u w=0.8u
m3702 70286 1837 VSS VSS nch l=0.04u w=0.8u
m3703 70287 1838 VSS VSS nch l=0.04u w=0.8u
m3704 70288 1839 VSS VSS nch l=0.04u w=0.8u
m3705 70289 1840 VSS VSS nch l=0.04u w=0.8u
m3706 70290 1841 VSS VSS nch l=0.04u w=0.8u
m3707 70291 1842 VSS VSS nch l=0.04u w=0.8u
m3708 70292 1843 VSS VSS nch l=0.04u w=0.8u
m3709 1875 FBDIV[5] 70278 VSS nch l=0.04u w=0.8u
m3710 1894 1934 VSS VSS nch l=0.04u w=0.4u
m3711 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3712 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3713 1876 1796 1860 VSS nch l=0.04u w=0.4u
m3714 1821 1983 70279 VSS nch l=0.04u w=0.8u
m3715 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3716 VSS 1909 70280 VSS nch l=0.04u w=0.12u
m3717 VSS 1910 70281 VSS nch l=0.04u w=0.12u
m3718 70293 11 1878 VSS nch l=0.04u w=0.8u
m3719 1899 3012 70282 VSS nch l=0.04u w=0.12u
m3720 1895 4328 1863 VSS nch l=0.04u w=0.4u
m3721 1896 4328 1864 VSS nch l=0.04u w=0.4u
m3722 1897 4328 1865 VSS nch l=0.04u w=0.4u
m3723 1898 4328 1866 VSS nch l=0.04u w=0.4u
m3724 1906 1854 VSS VSS nch l=0.04u w=0.4u
m3725 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3726 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3727 1900 4328 1868 VSS nch l=0.04u w=0.4u
m3728 1901 4328 1869 VSS nch l=0.04u w=0.4u
m3729 1902 4328 1870 VSS nch l=0.04u w=0.4u
m3730 70294 979 1879 VSS nch l=0.04u w=0.8u
m3731 1880 1720 70283 VSS nch l=0.04u w=0.8u
m3732 70295 1660 1881 VSS nch l=0.04u w=0.8u
m3733 1882 1722 70284 VSS nch l=0.04u w=0.8u
m3734 1903 4328 1872 VSS nch l=0.04u w=0.4u
m3735 1904 4328 1873 VSS nch l=0.04u w=0.4u
m3736 1905 4328 1874 VSS nch l=0.04u w=0.4u
m3737 70296 1657 1883 VSS nch l=0.04u w=0.8u
m3738 1884 1727 70285 VSS nch l=0.04u w=0.8u
m3739 1885 1728 70286 VSS nch l=0.04u w=0.8u
m3740 1886 1729 70287 VSS nch l=0.04u w=0.8u
m3741 70297 1577 1887 VSS nch l=0.04u w=0.8u
m3742 1888 1731 70288 VSS nch l=0.04u w=0.8u
m3743 1889 1732 70289 VSS nch l=0.04u w=0.8u
m3744 1890 1733 70290 VSS nch l=0.04u w=0.8u
m3745 70298 1579 1891 VSS nch l=0.04u w=0.8u
m3746 1892 1735 70291 VSS nch l=0.04u w=0.8u
m3747 1893 1736 70292 VSS nch l=0.04u w=0.8u
m3748 1908 94 VSS VSS nch l=0.04u w=0.4u
m3749 70299 1983 1821 VSS nch l=0.04u w=0.8u
m3750 1909 1861 VSS VSS nch l=0.04u w=0.4u
m3751 1910 1862 VSS VSS nch l=0.04u w=0.4u
m3752 VSS 1976 70293 VSS nch l=0.04u w=0.8u
m3753 1911 1917 1899 VSS nch l=0.04u w=0.4u
m3754 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3755 70300 1799 1895 VSS nch l=0.04u w=0.12u
m3756 70301 1800 1896 VSS nch l=0.04u w=0.12u
m3757 70302 1801 1897 VSS nch l=0.04u w=0.12u
m3758 70303 1802 1898 VSS nch l=0.04u w=0.12u
m3759 1912 1755 VSS VSS nch l=0.04u w=0.4u
m3760 70304 1807 1900 VSS nch l=0.04u w=0.12u
m3761 70305 1808 1901 VSS nch l=0.04u w=0.12u
m3762 70306 1809 1902 VSS nch l=0.04u w=0.12u
m3763 VSS 1657 70294 VSS nch l=0.04u w=0.8u
m3764 1913 1756 VSS VSS nch l=0.04u w=0.4u
m3765 VSS 139 70295 VSS nch l=0.04u w=0.8u
m3766 70307 1810 1903 VSS nch l=0.04u w=0.12u
m3767 70308 1811 1904 VSS nch l=0.04u w=0.12u
m3768 70309 1812 1905 VSS nch l=0.04u w=0.12u
m3769 VSS FRAC[19] 70296 VSS nch l=0.04u w=0.8u
m3770 VSS 1446 70297 VSS nch l=0.04u w=0.8u
m3771 VSS FRAC[19] 70298 VSS nch l=0.04u w=0.8u
m3772 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3773 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3774 70311 1850 VSS VSS nch l=0.04u w=0.8u
m3775 VSS 1934 1907 VSS nch l=0.04u w=0.4u
m3776 1915 377 VSS VSS nch l=0.04u w=0.4u
m3777 VSS 1936 70299 VSS nch l=0.04u w=0.8u
m3778 VSS 1679 VSS VSS nch l=0.26u w=0.8u
m3779 VSS 1941 70300 VSS nch l=0.04u w=0.12u
m3780 VSS 1505 70301 VSS nch l=0.04u w=0.12u
m3781 VSS 1942 70302 VSS nch l=0.04u w=0.12u
m3782 VSS 1508 70303 VSS nch l=0.04u w=0.12u
m3783 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3784 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3785 1918 1581 1912 VSS nch l=0.04u w=0.4u
m3786 VSS 688 70304 VSS nch l=0.04u w=0.12u
m3787 VSS 1789 70305 VSS nch l=0.04u w=0.12u
m3788 VSS 731 70306 VSS nch l=0.04u w=0.12u
m3789 458 1585 1913 VSS nch l=0.04u w=0.4u
m3790 VSS 1943 70307 VSS nch l=0.04u w=0.12u
m3791 VSS 1791 70308 VSS nch l=0.04u w=0.12u
m3792 VSS 735 70309 VSS nch l=0.04u w=0.12u
m3793 1920 1774 VSS VSS nch l=0.04u w=0.4u
m3794 1922 1776 VSS VSS nch l=0.04u w=0.4u
m3795 1924 1778 VSS VSS nch l=0.04u w=0.4u
m3796 1925 1780 VSS VSS nch l=0.04u w=0.4u
m3797 1926 1781 VSS VSS nch l=0.04u w=0.4u
m3798 1928 1783 VSS VSS nch l=0.04u w=0.4u
m3799 1929 1784 VSS VSS nch l=0.04u w=0.4u
m3800 1930 1785 VSS VSS nch l=0.04u w=0.4u
m3801 1932 1787 VSS VSS nch l=0.04u w=0.4u
m3802 1933 1788 VSS VSS nch l=0.04u w=0.4u
m3803 1914 1906 70311 VSS nch l=0.04u w=0.8u
m3804 1935 398 VSS VSS nch l=0.04u w=0.4u
m3805 1937 1938 VSS VSS nch l=0.04u w=0.8u
m3806 VSS 1694 VSS VSS nch l=0.26u w=0.8u
m3807 1939 4328 VSS VSS nch l=0.04u w=0.4u
m3808 1940 4328 VSS VSS nch l=0.04u w=0.4u
m3809 1941 1895 VSS VSS nch l=0.04u w=0.4u
m3810 1505 1896 VSS VSS nch l=0.04u w=0.4u
m3811 1942 1897 VSS VSS nch l=0.04u w=0.4u
m3812 1508 1898 VSS VSS nch l=0.04u w=0.4u
m3813 70318 303 1916 VSS nch l=0.04u w=0.8u
m3814 VSS 3012 1917 VSS nch l=0.04u w=0.4u
m3815 1581 1912 1918 VSS nch l=0.04u w=0.4u
m3816 688 1900 VSS VSS nch l=0.04u w=0.4u
m3817 1789 1901 VSS VSS nch l=0.04u w=0.4u
m3818 VSS 1704 VSS VSS nch l=0.26u w=0.8u
m3819 731 1902 VSS VSS nch l=0.04u w=0.4u
m3820 1585 1913 458 VSS nch l=0.04u w=0.4u
m3821 1943 1903 VSS VSS nch l=0.04u w=0.4u
m3822 1791 1904 VSS VSS nch l=0.04u w=0.4u
m3823 VSS 1706 VSS VSS nch l=0.26u w=0.8u
m3824 735 1905 VSS VSS nch l=0.04u w=0.4u
m3825 1820 1594 1920 VSS nch l=0.04u w=0.4u
m3826 1945 1595 1922 VSS nch l=0.04u w=0.4u
m3827 1790 1596 1924 VSS nch l=0.04u w=0.4u
m3828 1770 1597 1925 VSS nch l=0.04u w=0.4u
m3829 1947 1598 1926 VSS nch l=0.04u w=0.4u
m3830 1626 1599 1928 VSS nch l=0.04u w=0.4u
m3831 1805 1600 1929 VSS nch l=0.04u w=0.4u
m3832 1793 1601 1930 VSS nch l=0.04u w=0.4u
m3833 1628 1602 1932 VSS nch l=0.04u w=0.4u
m3834 1806 1603 1933 VSS nch l=0.04u w=0.4u
m3835 70320 1982 1934 VSS nch l=0.04u w=0.8u
m3836 70321 377 VSS VSS nch l=0.04u w=0.8u
m3837 70322 2079 1936 VSS nch l=0.04u w=0.8u
m3838 1952 1951 VSS VSS nch l=0.04u w=0.8u
m3839 VSS 149 70318 VSS nch l=0.04u w=0.8u
m3840 VSS 1714 VSS VSS nch l=0.26u w=0.8u
m3841 VSS 1717 VSS VSS nch l=0.26u w=0.8u
m3842 1953 1954 VSS VSS nch l=0.04u w=0.8u
m3843 1955 1956 VSS VSS nch l=0.04u w=0.8u
m3844 1594 1920 1820 VSS nch l=0.04u w=0.4u
m3845 1595 1922 1945 VSS nch l=0.04u w=0.4u
m3846 1596 1924 1790 VSS nch l=0.04u w=0.4u
m3847 1597 1925 1770 VSS nch l=0.04u w=0.4u
m3848 1598 1926 1947 VSS nch l=0.04u w=0.4u
m3849 1599 1928 1626 VSS nch l=0.04u w=0.4u
m3850 1600 1929 1805 VSS nch l=0.04u w=0.4u
m3851 1601 1930 1793 VSS nch l=0.04u w=0.4u
m3852 1602 1932 1628 VSS nch l=0.04u w=0.4u
m3853 1603 1933 1806 VSS nch l=0.04u w=0.4u
m3854 1819 1977 1919 VSS nch l=0.04u w=0.4u
m3855 1944 1978 1921 VSS nch l=0.04u w=0.4u
m3856 1946 1979 1923 VSS nch l=0.04u w=0.4u
m3857 1443 1980 1927 VSS nch l=0.04u w=0.4u
m3858 1445 1981 1931 VSS nch l=0.04u w=0.4u
m3859 70324 1914 VSS VSS nch l=0.04u w=0.8u
m3860 VSS 2648 70320 VSS nch l=0.04u w=0.8u
m3861 1948 REFDIV[3] 70321 VSS nch l=0.04u w=0.8u
m3862 VSS 2023 70322 VSS nch l=0.04u w=0.8u
m3863 1963 593 VSS VSS nch l=0.04u w=0.4u
m3864 VSS 1949 1949 VSS nch l=0.04u w=0.8u
m3865 1969 1968 VSS VSS nch l=0.04u w=0.8u
m3866 1970 1971 VSS VSS nch l=0.04u w=0.8u
m3867 1964 1939 1909 VSS nch l=0.04u w=0.4u
m3868 1965 1940 1910 VSS nch l=0.04u w=0.4u
m3869 1972 4328 VSS VSS nch l=0.04u w=0.4u
m3870 1973 4328 VSS VSS nch l=0.04u w=0.4u
m3871 1974 4328 VSS VSS nch l=0.04u w=0.4u
m3872 1975 4328 VSS VSS nch l=0.04u w=0.4u
m3873 70333 1593 1911 VSS nch l=0.04u w=0.8u
m3874 1977 1919 1819 VSS nch l=0.04u w=0.4u
m3875 1978 1921 1944 VSS nch l=0.04u w=0.4u
m3876 1979 1923 1946 VSS nch l=0.04u w=0.4u
m3877 1980 1927 1443 VSS nch l=0.04u w=0.4u
m3878 1981 1931 1445 VSS nch l=0.04u w=0.4u
m3879 1962 1875 70324 VSS nch l=0.04u w=0.8u
m3880 VSS 1967 1967 VSS nch l=0.04u w=0.8u
m3881 70351 4328 1964 VSS nch l=0.04u w=0.12u
m3882 70352 4328 1965 VSS nch l=0.04u w=0.12u
m3883 VSS 149 1976 VSS nch l=0.04u w=0.4u
m3884 VSS 1740 70333 VSS nch l=0.04u w=0.8u
m3885 70355 110 VSS VSS nch l=0.04u w=0.8u
m3886 VSS 1957 1977 VSS nch l=0.04u w=0.4u
m3887 70356 2022 VSS VSS nch l=0.04u w=0.8u
m3888 VSS 1958 1978 VSS nch l=0.04u w=0.4u
m3889 VSS 1959 1979 VSS nch l=0.04u w=0.4u
m3890 VSS 1960 1980 VSS nch l=0.04u w=0.4u
m3891 VSS 1961 1981 VSS nch l=0.04u w=0.4u
m3892 VSS 2021 1982 VSS nch l=0.04u w=0.4u
m3893 70357 1915 VSS VSS nch l=0.04u w=0.8u
m3894 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m3895 70358 REFDIV[4] 1983 VSS nch l=0.04u w=0.8u
m3896 1998 294 VSS VSS nch l=0.04u w=0.4u
m3897 VSS 2017 70351 VSS nch l=0.04u w=0.12u
m3898 VSS 2018 70352 VSS nch l=0.04u w=0.12u
m3899 VSS 1985 1985 VSS nch l=0.04u w=0.8u
m3900 VSS 1986 1986 VSS nch l=0.04u w=0.8u
m3901 1999 1972 1988 VSS nch l=0.04u w=0.4u
m3902 2000 1973 1947 VSS nch l=0.04u w=0.4u
m3903 2001 1974 1989 VSS nch l=0.04u w=0.4u
m3904 2002 1975 1793 VSS nch l=0.04u w=0.4u
m3905 1990 592 70355 VSS nch l=0.04u w=0.8u
m3906 1991 735 70356 VSS nch l=0.04u w=0.8u
m3907 VSS 1992 1992 VSS nch l=0.04u w=0.8u
m3908 70360 2073 VSS VSS nch l=0.04u w=0.8u
m3909 70361 2086 VSS VSS nch l=0.04u w=0.8u
m3910 70362 2616 VSS VSS nch l=0.04u w=0.8u
m3911 70363 2616 VSS VSS nch l=0.04u w=0.8u
m3912 VSS 1994 1994 VSS nch l=0.04u w=0.8u
m3913 70364 2616 VSS VSS nch l=0.04u w=0.8u
m3914 70365 FRAC[6] VSS VSS nch l=0.04u w=0.8u
m3915 VSS 2053 1996 VSS nch l=0.04u w=0.4u
m3916 70366 2074 VSS VSS nch l=0.04u w=0.8u
m3917 70367 2088 VSS VSS nch l=0.04u w=0.8u
m3918 70368 1989 VSS VSS nch l=0.04u w=0.8u
m3919 70369 1996 VSS VSS nch l=0.04u w=0.8u
m3920 70370 2089 VSS VSS nch l=0.04u w=0.8u
m3921 70371 FRAC[6] VSS VSS nch l=0.04u w=0.8u
m3922 70372 1996 VSS VSS nch l=0.04u w=0.8u
m3923 70373 1907 VSS VSS nch l=0.04u w=0.12u
m3924 1997 1860 70357 VSS nch l=0.04u w=0.8u
m3925 VSS 377 70358 VSS nch l=0.04u w=0.8u
m3926 110 2016 VSS VSS nch l=0.04u w=0.8u
m3927 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m3928 2017 1964 VSS VSS nch l=0.04u w=0.4u
m3929 2018 1965 VSS VSS nch l=0.04u w=0.4u
m3930 70374 4328 1999 VSS nch l=0.04u w=0.12u
m3931 70375 4328 2000 VSS nch l=0.04u w=0.12u
m3932 70376 4328 2001 VSS nch l=0.04u w=0.12u
m3933 70377 4328 2002 VSS nch l=0.04u w=0.12u
m3934 2019 3012 VSS VSS nch l=0.04u w=0.4u
m3935 2020 303 VSS VSS nch l=0.04u w=0.4u
m3936 70378 2158 1638 VSS nch l=0.04u w=0.8u
m3937 2003 2071 70360 VSS nch l=0.04u w=0.8u
m3938 70379 2160 1640 VSS nch l=0.04u w=0.8u
m3939 2004 2072 70361 VSS nch l=0.04u w=0.8u
m3940 2005 2223 70362 VSS nch l=0.04u w=0.8u
m3941 2006 2224 70363 VSS nch l=0.04u w=0.8u
m3942 2007 596 70364 VSS nch l=0.04u w=0.8u
m3943 70380 2162 1642 VSS nch l=0.04u w=0.8u
m3944 2008 2073 70365 VSS nch l=0.04u w=0.8u
m3945 2009 131 70366 VSS nch l=0.04u w=0.8u
m3946 2010 2074 70367 VSS nch l=0.04u w=0.8u
m3947 70381 2166 1646 VSS nch l=0.04u w=0.8u
m3948 2011 2075 70368 VSS nch l=0.04u w=0.8u
m3949 2012 2076 70369 VSS nch l=0.04u w=0.8u
m3950 2013 2077 70370 VSS nch l=0.04u w=0.8u
m3951 70382 2170 1650 VSS nch l=0.04u w=0.8u
m3952 2014 2078 70371 VSS nch l=0.04u w=0.8u
m3953 2015 FBDIV[6] 70372 VSS nch l=0.04u w=0.8u
m3954 2021 2151 70373 VSS nch l=0.04u w=0.12u
m3955 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m3956 2024 129 VSS VSS nch l=0.04u w=0.4u
m3957 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m3958 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m3959 VSS 2034 70374 VSS nch l=0.04u w=0.12u
m3960 VSS 2035 70375 VSS nch l=0.04u w=0.12u
m3961 VSS 2036 70376 VSS nch l=0.04u w=0.12u
m3962 VSS 2037 70377 VSS nch l=0.04u w=0.12u
m3963 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m3964 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m3965 2027 592 VSS VSS nch l=0.04u w=0.4u
m3966 VSS 2055 70378 VSS nch l=0.04u w=0.8u
m3967 2028 735 VSS VSS nch l=0.04u w=0.4u
m3968 VSS 2057 70379 VSS nch l=0.04u w=0.8u
m3969 VSS 2059 70380 VSS nch l=0.04u w=0.8u
m3970 VSS 2064 70381 VSS nch l=0.04u w=0.8u
m3971 VSS 2068 70382 VSS nch l=0.04u w=0.8u
m3972 2029 4328 VSS VSS nch l=0.04u w=0.4u
m3973 2030 2188 2021 VSS nch l=0.04u w=0.4u
m3974 VSS 3454 2022 VSS nch l=0.04u w=0.4u
m3975 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m3976 70386 1997 VSS VSS nch l=0.04u w=0.8u
m3977 VSS 377 2023 VSS nch l=0.04u w=0.4u
m3978 2032 4328 2017 VSS nch l=0.04u w=0.4u
m3979 2033 4328 2018 VSS nch l=0.04u w=0.4u
m3980 2034 1999 VSS VSS nch l=0.04u w=0.4u
m3981 2035 2000 VSS VSS nch l=0.04u w=0.4u
m3982 2036 2001 VSS VSS nch l=0.04u w=0.4u
m3983 2037 2002 VSS VSS nch l=0.04u w=0.4u
m3984 70387 2019 2025 VSS nch l=0.04u w=0.8u
m3985 70388 2020 2026 VSS nch l=0.04u w=0.8u
m3986 2038 110 2027 VSS nch l=0.04u w=0.4u
m3987 2039 2022 2028 VSS nch l=0.04u w=0.4u
m3988 2040 2071 VSS VSS nch l=0.04u w=0.4u
m3989 2041 2072 VSS VSS nch l=0.04u w=0.4u
m3990 2042 2005 VSS VSS nch l=0.04u w=0.4u
m3991 2043 2006 VSS VSS nch l=0.04u w=0.4u
m3992 2044 2007 VSS VSS nch l=0.04u w=0.4u
m3993 2045 2073 VSS VSS nch l=0.04u w=0.4u
m3994 2046 131 VSS VSS nch l=0.04u w=0.4u
m3995 2047 2074 VSS VSS nch l=0.04u w=0.4u
m3996 2048 2075 VSS VSS nch l=0.04u w=0.4u
m3997 2049 2076 VSS VSS nch l=0.04u w=0.4u
m3998 2050 2077 VSS VSS nch l=0.04u w=0.4u
m3999 2051 2078 VSS VSS nch l=0.04u w=0.4u
m4000 2052 FBDIV[6] VSS VSS nch l=0.04u w=0.4u
m4001 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m4002 2031 1948 70386 VSS nch l=0.04u w=0.8u
m4003 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m4004 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m4005 2054 441 VSS VSS nch l=0.04u w=0.4u
m4006 70389 1939 2032 VSS nch l=0.04u w=0.12u
m4007 70390 1940 2033 VSS nch l=0.04u w=0.12u
m4008 VSS 2270 70387 VSS nch l=0.04u w=0.8u
m4009 VSS 2271 70388 VSS nch l=0.04u w=0.8u
m4010 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m4011 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m4012 110 2027 2038 VSS nch l=0.04u w=0.4u
m4013 2022 2028 2039 VSS nch l=0.04u w=0.4u
m4014 70391 1919 VSS VSS nch l=0.04u w=0.8u
m4015 2056 2073 2040 VSS nch l=0.04u w=0.4u
m4016 70392 1921 VSS VSS nch l=0.04u w=0.8u
m4017 2058 2086 2041 VSS nch l=0.04u w=0.4u
m4018 70393 1923 VSS VSS nch l=0.04u w=0.8u
m4019 2060 FRAC[6] 2045 VSS nch l=0.04u w=0.4u
m4020 2062 2074 2046 VSS nch l=0.04u w=0.4u
m4021 2063 2088 2047 VSS nch l=0.04u w=0.4u
m4022 70394 1927 VSS VSS nch l=0.04u w=0.8u
m4023 2065 1989 2048 VSS nch l=0.04u w=0.4u
m4024 2066 1996 2049 VSS nch l=0.04u w=0.4u
m4025 2067 2089 2050 VSS nch l=0.04u w=0.4u
m4026 70395 1931 VSS VSS nch l=0.04u w=0.8u
m4027 2069 FRAC[6] 2051 VSS nch l=0.04u w=0.4u
m4028 2070 1996 2052 VSS nch l=0.04u w=0.4u
m4029 2061 2029 2053 VSS nch l=0.04u w=0.4u
m4030 70397 2122 2030 VSS nch l=0.04u w=0.8u
m4031 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m4032 70398 1948 2031 VSS nch l=0.04u w=0.8u
m4033 2079 2096 1677 VSS nch l=0.04u w=0.4u
m4034 VSS 60 70389 VSS nch l=0.04u w=0.12u
m4035 VSS 2098 70390 VSS nch l=0.04u w=0.12u
m4036 2080 4328 2034 VSS nch l=0.04u w=0.4u
m4037 2081 4328 2035 VSS nch l=0.04u w=0.4u
m4038 2082 4328 2036 VSS nch l=0.04u w=0.4u
m4039 2083 4328 2037 VSS nch l=0.04u w=0.4u
m4040 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m4041 2055 1957 70391 VSS nch l=0.04u w=0.8u
m4042 2073 2040 2056 VSS nch l=0.04u w=0.4u
m4043 2057 1958 70392 VSS nch l=0.04u w=0.8u
m4044 2086 2041 2058 VSS nch l=0.04u w=0.4u
m4045 2059 1959 70393 VSS nch l=0.04u w=0.8u
m4046 FRAC[6] 2045 2060 VSS nch l=0.04u w=0.4u
m4047 2074 2046 2062 VSS nch l=0.04u w=0.4u
m4048 2088 2047 2063 VSS nch l=0.04u w=0.4u
m4049 2064 1960 70394 VSS nch l=0.04u w=0.8u
m4050 1989 2048 2065 VSS nch l=0.04u w=0.4u
m4051 1996 2049 2066 VSS nch l=0.04u w=0.4u
m4052 2089 2050 2067 VSS nch l=0.04u w=0.4u
m4053 2068 1961 70395 VSS nch l=0.04u w=0.8u
m4054 FRAC[6] 2051 2069 VSS nch l=0.04u w=0.4u
m4055 1996 2052 2070 VSS nch l=0.04u w=0.4u
m4056 2090 4328 VSS VSS nch l=0.04u w=0.4u
m4057 2091 4328 VSS VSS nch l=0.04u w=0.4u
m4058 2092 4328 VSS VSS nch l=0.04u w=0.4u
m4059 2093 4328 VSS VSS nch l=0.04u w=0.4u
m4060 2094 4328 VSS VSS nch l=0.04u w=0.4u
m4061 2095 4328 VSS VSS nch l=0.04u w=0.4u
m4062 70399 4328 2061 VSS nch l=0.04u w=0.12u
m4063 VSS 2648 70397 VSS nch l=0.04u w=0.8u
m4064 VSS 1997 70398 VSS nch l=0.04u w=0.8u
m4065 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m4066 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m4067 2096 1677 2079 VSS nch l=0.04u w=0.4u
m4068 2097 735 VSS VSS nch l=0.04u w=0.4u
m4069 60 2032 VSS VSS nch l=0.04u w=0.4u
m4070 2098 2033 VSS VSS nch l=0.04u w=0.4u
m4071 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m4072 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m4073 70403 1972 2080 VSS nch l=0.04u w=0.12u
m4074 70404 1973 2081 VSS nch l=0.04u w=0.12u
m4075 70405 1974 2082 VSS nch l=0.04u w=0.12u
m4076 70406 1975 2083 VSS nch l=0.04u w=0.12u
m4077 VSS 4353 2084 VSS nch l=0.04u w=0.4u
m4078 VSS 11 2085 VSS nch l=0.04u w=0.4u
m4079 VSS 2111 70399 VSS nch l=0.04u w=0.12u
m4080 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m4081 70407 2030 VSS VSS nch l=0.04u w=0.24u
m4082 VSS 2075 70403 VSS nch l=0.04u w=0.12u
m4083 VSS 1792 70404 VSS nch l=0.04u w=0.12u
m4084 VSS 2078 70405 VSS nch l=0.04u w=0.12u
m4085 VSS 1794 70406 VSS nch l=0.04u w=0.12u
m4086 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m4087 70423 2038 2099 VSS nch l=0.04u w=0.8u
m4088 70424 2039 2100 VSS nch l=0.04u w=0.8u
m4089 2111 2061 VSS VSS nch l=0.04u w=0.4u
m4090 2122 2188 70407 VSS nch l=0.04u w=0.24u
m4091 2105 2090 2102 VSS nch l=0.04u w=0.4u
m4092 2106 2091 2103 VSS nch l=0.04u w=0.4u
m4093 2107 2092 595 VSS nch l=0.04u w=0.4u
m4094 2108 2093 2042 VSS nch l=0.04u w=0.4u
m4095 2109 2094 2043 VSS nch l=0.04u w=0.4u
m4096 2110 2095 2044 VSS nch l=0.04u w=0.4u
m4097 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m4098 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m4099 2123 76 VSS VSS nch l=0.04u w=0.4u
m4100 VSS 2096 2104 VSS nch l=0.04u w=0.4u
m4101 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m4102 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m4103 139 1027 VSS VSS nch l=0.04u w=0.4u
m4104 2124 2131 VSS VSS nch l=0.04u w=0.4u
m4105 2125 1099 VSS VSS nch l=0.04u w=0.4u
m4106 2075 2080 VSS VSS nch l=0.04u w=0.4u
m4107 1792 2081 VSS VSS nch l=0.04u w=0.4u
m4108 2078 2082 VSS VSS nch l=0.04u w=0.4u
m4109 1794 2083 VSS VSS nch l=0.04u w=0.4u
m4110 2126 2084 2025 VSS nch l=0.04u w=0.4u
m4111 2127 2085 2026 VSS nch l=0.04u w=0.4u
m4112 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m4113 VSS 1867 70423 VSS nch l=0.04u w=0.8u
m4114 VSS 1871 70424 VSS nch l=0.04u w=0.8u
m4115 1934 2151 2122 VSS nch l=0.04u w=0.4u
m4116 70425 4328 2105 VSS nch l=0.04u w=0.12u
m4117 70426 4328 2106 VSS nch l=0.04u w=0.12u
m4118 70427 4328 2107 VSS nch l=0.04u w=0.12u
m4119 1957 2133 1943 VSS nch l=0.04u w=0.4u
m4120 70428 2056 2112 VSS nch l=0.04u w=0.8u
m4121 1958 2134 139 VSS nch l=0.04u w=0.4u
m4122 70429 2058 2113 VSS nch l=0.04u w=0.8u
m4123 70430 4328 2108 VSS nch l=0.04u w=0.12u
m4124 70431 4328 2109 VSS nch l=0.04u w=0.12u
m4125 70432 4328 2110 VSS nch l=0.04u w=0.12u
m4126 1959 2135 FRAC[18] VSS nch l=0.04u w=0.4u
m4127 70433 2060 2114 VSS nch l=0.04u w=0.8u
m4128 70434 2062 2115 VSS nch l=0.04u w=0.8u
m4129 70435 2063 2116 VSS nch l=0.04u w=0.8u
m4130 1960 2136 1445 VSS nch l=0.04u w=0.4u
m4131 70436 2065 2117 VSS nch l=0.04u w=0.8u
m4132 70437 2066 2118 VSS nch l=0.04u w=0.8u
m4133 70438 2067 2119 VSS nch l=0.04u w=0.8u
m4134 1961 2137 FRAC[18] VSS nch l=0.04u w=0.4u
m4135 70439 2069 2120 VSS nch l=0.04u w=0.8u
m4136 70440 2070 2121 VSS nch l=0.04u w=0.8u
m4137 2128 155 VSS VSS nch l=0.04u w=0.4u
m4138 2129 60 2124 VSS nch l=0.04u w=0.4u
m4139 2130 2098 2125 VSS nch l=0.04u w=0.4u
m4140 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m4141 70441 4353 2126 VSS nch l=0.04u w=0.24u
m4142 70442 11 2127 VSS nch l=0.04u w=0.24u
m4143 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m4144 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m4145 VSS 2144 70425 VSS nch l=0.04u w=0.12u
m4146 VSS 2145 70426 VSS nch l=0.04u w=0.12u
m4147 VSS 2146 70427 VSS nch l=0.04u w=0.12u
m4148 2133 1943 1957 VSS nch l=0.04u w=0.4u
m4149 VSS 1880 70428 VSS nch l=0.04u w=0.8u
m4150 2134 139 1958 VSS nch l=0.04u w=0.4u
m4151 VSS 1882 70429 VSS nch l=0.04u w=0.8u
m4152 VSS 2148 70430 VSS nch l=0.04u w=0.12u
m4153 VSS 2149 70431 VSS nch l=0.04u w=0.12u
m4154 VSS 2150 70432 VSS nch l=0.04u w=0.12u
m4155 2135 FRAC[18] 1959 VSS nch l=0.04u w=0.4u
m4156 VSS 1884 70433 VSS nch l=0.04u w=0.8u
m4157 2132 4328 2111 VSS nch l=0.04u w=0.4u
m4158 VSS 1885 70434 VSS nch l=0.04u w=0.8u
m4159 VSS 1886 70435 VSS nch l=0.04u w=0.8u
m4160 2136 1445 1960 VSS nch l=0.04u w=0.4u
m4161 VSS 1888 70436 VSS nch l=0.04u w=0.8u
m4162 VSS 1889 70437 VSS nch l=0.04u w=0.8u
m4163 VSS 1890 70438 VSS nch l=0.04u w=0.8u
m4164 2137 FRAC[18] 1961 VSS nch l=0.04u w=0.4u
m4165 VSS 1892 70439 VSS nch l=0.04u w=0.8u
m4166 VSS 1893 70440 VSS nch l=0.04u w=0.8u
m4167 2138 2123 2031 VSS nch l=0.04u w=0.4u
m4168 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m4169 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m4170 70443 683 2096 VSS nch l=0.04u w=0.8u
m4171 60 2124 2129 VSS nch l=0.04u w=0.4u
m4172 2098 2125 2130 VSS nch l=0.04u w=0.4u
m4173 140 3338 VSS VSS nch l=0.04u w=0.4u
m4174 2139 4328 VSS VSS nch l=0.04u w=0.4u
m4175 2140 4328 VSS VSS nch l=0.04u w=0.4u
m4176 2141 4328 VSS VSS nch l=0.04u w=0.4u
m4177 2142 4328 VSS VSS nch l=0.04u w=0.4u
m4178 VSS 2156 70441 VSS nch l=0.04u w=0.24u
m4179 VSS 2157 70442 VSS nch l=0.04u w=0.24u
m4180 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m4181 70444 2099 VSS VSS nch l=0.04u w=0.8u
m4182 2144 2105 VSS VSS nch l=0.04u w=0.4u
m4183 2145 2106 VSS VSS nch l=0.04u w=0.4u
m4184 2146 2107 VSS VSS nch l=0.04u w=0.4u
m4185 VSS 688 2133 VSS nch l=0.04u w=0.4u
m4186 70445 2100 VSS VSS nch l=0.04u w=0.8u
m4187 VSS 1946 2134 VSS nch l=0.04u w=0.4u
m4188 2148 2108 VSS VSS nch l=0.04u w=0.4u
m4189 2149 2109 VSS VSS nch l=0.04u w=0.4u
m4190 2150 2110 VSS VSS nch l=0.04u w=0.4u
m4191 VSS 1943 2135 VSS nch l=0.04u w=0.4u
m4192 70446 2029 2132 VSS nch l=0.04u w=0.12u
m4193 VSS 1576 2136 VSS nch l=0.04u w=0.4u
m4194 VSS 1578 2137 VSS nch l=0.04u w=0.4u
m4195 2151 2188 VSS VSS nch l=0.04u w=0.4u
m4196 70447 155 VSS VSS nch l=0.04u w=0.8u
m4197 70448 76 2138 VSS nch l=0.04u w=0.12u
m4198 70449 1240 70443 VSS nch l=0.04u w=0.8u
m4199 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m4200 70450 2716 VSS VSS nch l=0.04u w=0.8u
m4201 70451 2716 VSS VSS nch l=0.04u w=0.8u
m4202 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m4203 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m4204 2143 1990 70444 VSS nch l=0.04u w=0.8u
m4205 2147 1991 70445 VSS nch l=0.04u w=0.8u
m4206 VSS 2184 70446 VSS nch l=0.04u w=0.12u
m4207 70452 2112 VSS VSS nch l=0.04u w=0.8u
m4208 70453 2113 VSS VSS nch l=0.04u w=0.8u
m4209 70454 2114 VSS VSS nch l=0.04u w=0.8u
m4210 70455 2115 VSS VSS nch l=0.04u w=0.8u
m4211 70456 2116 VSS VSS nch l=0.04u w=0.8u
m4212 70457 2117 VSS VSS nch l=0.04u w=0.8u
m4213 70458 2118 VSS VSS nch l=0.04u w=0.8u
m4214 70459 2119 VSS VSS nch l=0.04u w=0.8u
m4215 70460 2120 VSS VSS nch l=0.04u w=0.8u
m4216 70461 2121 VSS VSS nch l=0.04u w=0.8u
m4217 2152 FBDIV[6] 70447 VSS nch l=0.04u w=0.8u
m4218 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m4219 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m4220 VSS 2185 70448 VSS nch l=0.04u w=0.12u
m4221 VSS 2194 70449 VSS nch l=0.04u w=0.8u
m4222 459 3610 VSS VSS nch l=0.04u w=0.4u
m4223 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m4224 2174 2139 2153 VSS nch l=0.04u w=0.4u
m4225 2175 2140 2154 VSS nch l=0.04u w=0.4u
m4226 2176 2141 2155 VSS nch l=0.04u w=0.4u
m4227 2177 2142 2076 VSS nch l=0.04u w=0.4u
m4228 2156 2126 70450 VSS nch l=0.04u w=0.8u
m4229 2157 2127 70451 VSS nch l=0.04u w=0.8u
m4230 2184 2132 VSS VSS nch l=0.04u w=0.4u
m4231 2178 4328 2144 VSS nch l=0.04u w=0.4u
m4232 2179 4328 2145 VSS nch l=0.04u w=0.4u
m4233 2180 4328 2146 VSS nch l=0.04u w=0.4u
m4234 70462 688 2158 VSS nch l=0.04u w=0.8u
m4235 2159 2003 70452 VSS nch l=0.04u w=0.8u
m4236 70463 1946 2160 VSS nch l=0.04u w=0.8u
m4237 2161 2004 70453 VSS nch l=0.04u w=0.8u
m4238 2181 4328 2148 VSS nch l=0.04u w=0.4u
m4239 2182 4328 2149 VSS nch l=0.04u w=0.4u
m4240 2183 4328 2150 VSS nch l=0.04u w=0.4u
m4241 70464 1943 2162 VSS nch l=0.04u w=0.8u
m4242 2163 2008 70454 VSS nch l=0.04u w=0.8u
m4243 2164 2009 70455 VSS nch l=0.04u w=0.8u
m4244 2165 2010 70456 VSS nch l=0.04u w=0.8u
m4245 70465 1576 2166 VSS nch l=0.04u w=0.8u
m4246 2167 2011 70457 VSS nch l=0.04u w=0.8u
m4247 2168 2012 70458 VSS nch l=0.04u w=0.8u
m4248 2169 2013 70459 VSS nch l=0.04u w=0.8u
m4249 70466 1578 2170 VSS nch l=0.04u w=0.8u
m4250 2171 2014 70460 VSS nch l=0.04u w=0.8u
m4251 2172 2015 70461 VSS nch l=0.04u w=0.8u
m4252 VSS 2188 2173 VSS nch l=0.04u w=0.4u
m4253 2185 2138 VSS VSS nch l=0.04u w=0.4u
m4254 VSS 1950 VSS VSS nch l=0.26u w=0.8u
m4255 70467 4328 2174 VSS nch l=0.04u w=0.12u
m4256 70468 4328 2175 VSS nch l=0.04u w=0.12u
m4257 70469 4328 2176 VSS nch l=0.04u w=0.12u
m4258 70470 4328 2177 VSS nch l=0.04u w=0.12u
m4259 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m4260 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m4261 2186 2038 VSS VSS nch l=0.04u w=0.4u
m4262 70471 2090 2178 VSS nch l=0.04u w=0.12u
m4263 70472 2091 2179 VSS nch l=0.04u w=0.12u
m4264 70473 2092 2180 VSS nch l=0.04u w=0.12u
m4265 VSS 1943 70462 VSS nch l=0.04u w=0.8u
m4266 2187 2039 VSS VSS nch l=0.04u w=0.4u
m4267 VSS 139 70463 VSS nch l=0.04u w=0.8u
m4268 70474 2093 2181 VSS nch l=0.04u w=0.12u
m4269 70475 2094 2182 VSS nch l=0.04u w=0.12u
m4270 70476 2095 2183 VSS nch l=0.04u w=0.12u
m4271 VSS FRAC[18] 70464 VSS nch l=0.04u w=0.8u
m4272 VSS 1445 70465 VSS nch l=0.04u w=0.8u
m4273 VSS FRAC[18] 70466 VSS nch l=0.04u w=0.8u
m4274 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m4275 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m4276 70478 2128 VSS VSS nch l=0.04u w=0.8u
m4277 2190 2191 VSS VSS nch l=0.04u w=0.8u
m4278 2192 4328 VSS VSS nch l=0.04u w=0.4u
m4279 2193 4328 VSS VSS nch l=0.04u w=0.4u
m4280 2194 2228 VSS VSS nch l=0.04u w=0.4u
m4281 VSS 1966 VSS VSS nch l=0.26u w=0.8u
m4282 VSS 2218 70467 VSS nch l=0.04u w=0.12u
m4283 VSS 2219 70468 VSS nch l=0.04u w=0.12u
m4284 VSS 2220 70469 VSS nch l=0.04u w=0.12u
m4285 VSS 2221 70470 VSS nch l=0.04u w=0.12u
m4286 755 3760 VSS VSS nch l=0.04u w=0.4u
m4287 2195 4353 2156 VSS nch l=0.04u w=0.4u
m4288 2196 11 2157 VSS nch l=0.04u w=0.4u
m4289 2197 1867 2186 VSS nch l=0.04u w=0.4u
m4290 VSS 395 70471 VSS nch l=0.04u w=0.12u
m4291 VSS 2071 70472 VSS nch l=0.04u w=0.12u
m4292 VSS 437 70473 VSS nch l=0.04u w=0.12u
m4293 754 1871 2187 VSS nch l=0.04u w=0.4u
m4294 VSS 2222 70474 VSS nch l=0.04u w=0.12u
m4295 VSS 2073 70475 VSS nch l=0.04u w=0.12u
m4296 VSS 441 70476 VSS nch l=0.04u w=0.12u
m4297 2199 2056 VSS VSS nch l=0.04u w=0.4u
m4298 2201 2058 VSS VSS nch l=0.04u w=0.4u
m4299 2203 2060 VSS VSS nch l=0.04u w=0.4u
m4300 2204 2062 VSS VSS nch l=0.04u w=0.4u
m4301 2205 2063 VSS VSS nch l=0.04u w=0.4u
m4302 2207 2065 VSS VSS nch l=0.04u w=0.4u
m4303 2208 2066 VSS VSS nch l=0.04u w=0.4u
m4304 2209 2067 VSS VSS nch l=0.04u w=0.4u
m4305 2211 2069 VSS VSS nch l=0.04u w=0.4u
m4306 2212 2070 VSS VSS nch l=0.04u w=0.4u
m4307 70480 2244 2188 VSS nch l=0.04u w=0.8u
m4308 2189 2184 70478 VSS nch l=0.04u w=0.8u
m4309 2213 76 2185 VSS nch l=0.04u w=0.4u
m4310 VSS 2228 2194 VSS nch l=0.04u w=0.4u
m4311 2217 2216 VSS VSS nch l=0.04u w=0.8u
m4312 2218 2174 VSS VSS nch l=0.04u w=0.4u
m4313 2219 2175 VSS VSS nch l=0.04u w=0.4u
m4314 2220 2176 VSS VSS nch l=0.04u w=0.4u
m4315 2221 2177 VSS VSS nch l=0.04u w=0.4u
m4316 VSS 1984 VSS VSS nch l=0.26u w=0.8u
m4317 VSS 1987 VSS VSS nch l=0.26u w=0.8u
m4318 70486 2084 2195 VSS nch l=0.04u w=0.12u
m4319 70487 2085 2196 VSS nch l=0.04u w=0.12u
m4320 1867 2186 2197 VSS nch l=0.04u w=0.4u
m4321 395 2178 VSS VSS nch l=0.04u w=0.4u
m4322 2071 2179 VSS VSS nch l=0.04u w=0.4u
m4323 VSS 1993 VSS VSS nch l=0.26u w=0.8u
m4324 437 2180 VSS VSS nch l=0.04u w=0.4u
m4325 1871 2187 754 VSS nch l=0.04u w=0.4u
m4326 2222 2181 VSS VSS nch l=0.04u w=0.4u
m4327 2073 2182 VSS VSS nch l=0.04u w=0.4u
m4328 VSS 1995 VSS VSS nch l=0.26u w=0.8u
m4329 441 2183 VSS VSS nch l=0.04u w=0.4u
m4330 2103 1880 2199 VSS nch l=0.04u w=0.4u
m4331 2224 1882 2201 VSS nch l=0.04u w=0.4u
m4332 2072 1884 2203 VSS nch l=0.04u w=0.4u
m4333 2053 1885 2204 VSS nch l=0.04u w=0.4u
m4334 2154 1886 2205 VSS nch l=0.04u w=0.4u
m4335 1988 1888 2207 VSS nch l=0.04u w=0.4u
m4336 2088 1889 2208 VSS nch l=0.04u w=0.4u
m4337 2076 1890 2209 VSS nch l=0.04u w=0.4u
m4338 1989 1892 2211 VSS nch l=0.04u w=0.4u
m4339 2089 1893 2212 VSS nch l=0.04u w=0.4u
m4340 VSS 2648 70480 VSS nch l=0.04u w=0.8u
m4341 70489 2123 2213 VSS nch l=0.04u w=0.12u
m4342 VSS 2214 2214 VSS nch l=0.04u w=0.8u
m4343 2226 2192 2129 VSS nch l=0.04u w=0.4u
m4344 2227 2193 2130 VSS nch l=0.04u w=0.4u
m4345 2232 2231 VSS VSS nch l=0.04u w=0.8u
m4346 2233 2234 VSS VSS nch l=0.04u w=0.8u
m4347 VSS 2300 70486 VSS nch l=0.04u w=0.12u
m4348 VSS 2301 70487 VSS nch l=0.04u w=0.12u
m4349 1042 3479 VSS VSS nch l=0.04u w=0.4u
m4350 2235 2236 VSS VSS nch l=0.04u w=0.8u
m4351 2237 2238 VSS VSS nch l=0.04u w=0.8u
m4352 1880 2199 2103 VSS nch l=0.04u w=0.4u
m4353 1882 2201 2224 VSS nch l=0.04u w=0.4u
m4354 1884 2203 2072 VSS nch l=0.04u w=0.4u
m4355 1885 2204 2053 VSS nch l=0.04u w=0.4u
m4356 1886 2205 2154 VSS nch l=0.04u w=0.4u
m4357 1888 2207 1988 VSS nch l=0.04u w=0.4u
m4358 1889 2208 2088 VSS nch l=0.04u w=0.4u
m4359 1890 2209 2076 VSS nch l=0.04u w=0.4u
m4360 1892 2211 1989 VSS nch l=0.04u w=0.4u
m4361 1893 2212 2089 VSS nch l=0.04u w=0.4u
m4362 2102 2256 2198 VSS nch l=0.04u w=0.4u
m4363 2223 2257 2200 VSS nch l=0.04u w=0.4u
m4364 2225 2258 2202 VSS nch l=0.04u w=0.4u
m4365 1814 2259 2206 VSS nch l=0.04u w=0.4u
m4366 1815 2260 2210 VSS nch l=0.04u w=0.4u
m4367 70491 2189 VSS VSS nch l=0.04u w=0.8u
m4368 VSS 1876 70489 VSS nch l=0.04u w=0.12u
m4369 70500 4328 2226 VSS nch l=0.04u w=0.12u
m4370 70501 4328 2227 VSS nch l=0.04u w=0.12u
m4371 70502 1742 2228 VSS nch l=0.04u w=0.8u
m4372 VSS 2230 2230 VSS nch l=0.04u w=0.8u
m4373 2246 4328 2218 VSS nch l=0.04u w=0.4u
m4374 2247 4328 2219 VSS nch l=0.04u w=0.4u
m4375 2248 4328 2220 VSS nch l=0.04u w=0.4u
m4376 2249 4328 2221 VSS nch l=0.04u w=0.4u
m4377 2250 2195 VSS VSS nch l=0.04u w=0.4u
m4378 2251 2196 VSS VSS nch l=0.04u w=0.4u
m4379 2256 2198 2102 VSS nch l=0.04u w=0.4u
m4380 2257 2200 2223 VSS nch l=0.04u w=0.4u
m4381 2258 2202 2225 VSS nch l=0.04u w=0.4u
m4382 2259 2206 1814 VSS nch l=0.04u w=0.4u
m4383 2260 2210 1815 VSS nch l=0.04u w=0.4u
m4384 VSS 2285 2244 VSS nch l=0.04u w=0.4u
m4385 2245 2152 70491 VSS nch l=0.04u w=0.8u
m4386 1876 2213 VSS VSS nch l=0.04u w=0.4u
m4387 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4388 VSS 2268 70500 VSS nch l=0.04u w=0.12u
m4389 VSS 2269 70501 VSS nch l=0.04u w=0.12u
m4390 VSS 2286 70502 VSS nch l=0.04u w=0.8u
m4391 70519 2139 2246 VSS nch l=0.04u w=0.12u
m4392 70520 2140 2247 VSS nch l=0.04u w=0.12u
m4393 70521 2141 2248 VSS nch l=0.04u w=0.12u
m4394 70522 2142 2249 VSS nch l=0.04u w=0.12u
m4395 VSS 2253 2253 VSS nch l=0.04u w=0.8u
m4396 VSS 2254 2254 VSS nch l=0.04u w=0.8u
m4397 1514 3204 VSS VSS nch l=0.04u w=0.4u
m4398 70526 110 VSS VSS nch l=0.04u w=0.8u
m4399 VSS 2239 2256 VSS nch l=0.04u w=0.4u
m4400 70527 2290 VSS VSS nch l=0.04u w=0.8u
m4401 VSS 2240 2257 VSS nch l=0.04u w=0.4u
m4402 VSS 2241 2258 VSS nch l=0.04u w=0.4u
m4403 VSS 2242 2259 VSS nch l=0.04u w=0.4u
m4404 VSS 2243 2260 VSS nch l=0.04u w=0.4u
m4405 70528 2173 VSS VSS nch l=0.04u w=0.12u
m4406 2268 2226 VSS VSS nch l=0.04u w=0.4u
m4407 2269 2227 VSS VSS nch l=0.04u w=0.4u
m4408 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4409 VSS 2287 70519 VSS nch l=0.04u w=0.12u
m4410 VSS 2074 70520 VSS nch l=0.04u w=0.12u
m4411 VSS 2288 70521 VSS nch l=0.04u w=0.12u
m4412 VSS 2077 70522 VSS nch l=0.04u w=0.12u
m4413 70529 2716 VSS VSS nch l=0.04u w=0.8u
m4414 70530 2716 VSS VSS nch l=0.04u w=0.8u
m4415 2261 292 70526 VSS nch l=0.04u w=0.8u
m4416 2262 1027 70527 VSS nch l=0.04u w=0.8u
m4417 2285 2403 70528 VSS nch l=0.04u w=0.12u
m4418 VSS 2263 2263 VSS nch l=0.04u w=0.8u
m4419 70533 2344 VSS VSS nch l=0.04u w=0.8u
m4420 70534 2357 VSS VSS nch l=0.04u w=0.8u
m4421 70535 2616 VSS VSS nch l=0.04u w=0.8u
m4422 70536 2616 VSS VSS nch l=0.04u w=0.8u
m4423 VSS 2265 2265 VSS nch l=0.04u w=0.8u
m4424 70537 2616 VSS VSS nch l=0.04u w=0.8u
m4425 70538 FRAC[7] VSS VSS nch l=0.04u w=0.8u
m4426 VSS 2321 2267 VSS nch l=0.04u w=0.4u
m4427 70539 2345 VSS VSS nch l=0.04u w=0.8u
m4428 70540 2359 VSS VSS nch l=0.04u w=0.8u
m4429 70541 2324 VSS VSS nch l=0.04u w=0.8u
m4430 70542 2267 VSS VSS nch l=0.04u w=0.8u
m4431 70543 2360 VSS VSS nch l=0.04u w=0.8u
m4432 70544 FRAC[7] VSS VSS nch l=0.04u w=0.8u
m4433 70545 2267 VSS VSS nch l=0.04u w=0.8u
m4434 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4435 2286 1876 VSS VSS nch l=0.04u w=0.4u
m4436 VSS 2252 VSS VSS nch l=0.26u w=0.8u
m4437 VSS 2255 VSS VSS nch l=0.26u w=0.8u
m4438 2287 2246 VSS VSS nch l=0.04u w=0.4u
m4439 2074 2247 VSS VSS nch l=0.04u w=0.4u
m4440 2288 2248 VSS VSS nch l=0.04u w=0.4u
m4441 2077 2249 VSS VSS nch l=0.04u w=0.4u
m4442 2270 2250 70529 VSS nch l=0.04u w=0.8u
m4443 2271 2251 70530 VSS nch l=0.04u w=0.8u
m4444 1803 2925 VSS VSS nch l=0.04u w=0.4u
m4445 2289 2454 2285 VSS nch l=0.04u w=0.4u
m4446 70547 2428 1919 VSS nch l=0.04u w=0.8u
m4447 2272 2342 70533 VSS nch l=0.04u w=0.8u
m4448 70548 2430 1921 VSS nch l=0.04u w=0.8u
m4449 2273 2343 70534 VSS nch l=0.04u w=0.8u
m4450 2274 2488 70535 VSS nch l=0.04u w=0.8u
m4451 2275 2489 70536 VSS nch l=0.04u w=0.8u
m4452 2276 297 70537 VSS nch l=0.04u w=0.8u
m4453 70549 2432 1923 VSS nch l=0.04u w=0.8u
m4454 2277 2344 70538 VSS nch l=0.04u w=0.8u
m4455 2278 131 70539 VSS nch l=0.04u w=0.8u
m4456 2279 2345 70540 VSS nch l=0.04u w=0.8u
m4457 70550 2436 1927 VSS nch l=0.04u w=0.8u
m4458 2280 2346 70541 VSS nch l=0.04u w=0.8u
m4459 2281 2325 70542 VSS nch l=0.04u w=0.8u
m4460 2282 2347 70543 VSS nch l=0.04u w=0.8u
m4461 70551 2440 1931 VSS nch l=0.04u w=0.8u
m4462 2283 2348 70544 VSS nch l=0.04u w=0.8u
m4463 2284 FBDIV[7] 70545 VSS nch l=0.04u w=0.8u
m4464 VSS 1876 2286 VSS nch l=0.04u w=0.4u
m4465 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4466 2291 4328 2268 VSS nch l=0.04u w=0.4u
m4467 2292 4328 2269 VSS nch l=0.04u w=0.4u
m4468 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4469 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4470 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4471 2293 292 VSS VSS nch l=0.04u w=0.4u
m4472 VSS 2326 70547 VSS nch l=0.04u w=0.8u
m4473 2294 1027 VSS VSS nch l=0.04u w=0.4u
m4474 VSS 2328 70548 VSS nch l=0.04u w=0.8u
m4475 VSS 2330 70549 VSS nch l=0.04u w=0.8u
m4476 VSS 2335 70550 VSS nch l=0.04u w=0.8u
m4477 VSS 2339 70551 VSS nch l=0.04u w=0.8u
m4478 2295 4328 VSS VSS nch l=0.04u w=0.4u
m4479 VSS 3736 2290 VSS nch l=0.04u w=0.4u
m4480 VSS 2252 VSS VSS nch l=0.26u w=0.8u
m4481 VSS 2255 VSS VSS nch l=0.26u w=0.8u
m4482 70557 2192 2291 VSS nch l=0.04u w=0.12u
m4483 70558 2193 2292 VSS nch l=0.04u w=0.12u
m4484 2296 4328 VSS VSS nch l=0.04u w=0.4u
m4485 2297 4328 VSS VSS nch l=0.04u w=0.4u
m4486 2298 4328 VSS VSS nch l=0.04u w=0.4u
m4487 2299 4328 VSS VSS nch l=0.04u w=0.4u
m4488 2300 2270 VSS VSS nch l=0.04u w=0.4u
m4489 2301 2271 VSS VSS nch l=0.04u w=0.4u
m4490 2086 2486 VSS VSS nch l=0.04u w=0.4u
m4491 2302 110 2293 VSS nch l=0.04u w=0.4u
m4492 2303 2290 2294 VSS nch l=0.04u w=0.4u
m4493 70559 2369 2289 VSS nch l=0.04u w=0.8u
m4494 2308 2342 VSS VSS nch l=0.04u w=0.4u
m4495 2309 2343 VSS VSS nch l=0.04u w=0.4u
m4496 2310 2274 VSS VSS nch l=0.04u w=0.4u
m4497 2311 2275 VSS VSS nch l=0.04u w=0.4u
m4498 2312 2276 VSS VSS nch l=0.04u w=0.4u
m4499 2313 2344 VSS VSS nch l=0.04u w=0.4u
m4500 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4501 2314 131 VSS VSS nch l=0.04u w=0.4u
m4502 2315 2345 VSS VSS nch l=0.04u w=0.4u
m4503 2316 2346 VSS VSS nch l=0.04u w=0.4u
m4504 2317 2325 VSS VSS nch l=0.04u w=0.4u
m4505 2318 2347 VSS VSS nch l=0.04u w=0.4u
m4506 2319 2348 VSS VSS nch l=0.04u w=0.4u
m4507 2320 FBDIV[7] VSS VSS nch l=0.04u w=0.4u
m4508 VSS 2349 70557 VSS nch l=0.04u w=0.12u
m4509 VSS 2350 70558 VSS nch l=0.04u w=0.12u
m4510 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4511 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4512 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4513 110 2293 2302 VSS nch l=0.04u w=0.4u
m4514 2290 2294 2303 VSS nch l=0.04u w=0.4u
m4515 VSS 2304 2304 VSS nch l=0.04u w=0.8u
m4516 VSS 2307 2307 VSS nch l=0.04u w=0.8u
m4517 VSS 2648 70559 VSS nch l=0.04u w=0.8u
m4518 70560 2198 VSS VSS nch l=0.04u w=0.8u
m4519 2327 2344 2308 VSS nch l=0.04u w=0.4u
m4520 70561 2200 VSS VSS nch l=0.04u w=0.8u
m4521 2329 2357 2309 VSS nch l=0.04u w=0.4u
m4522 70562 2202 VSS VSS nch l=0.04u w=0.8u
m4523 2331 FRAC[7] 2313 VSS nch l=0.04u w=0.4u
m4524 2333 2345 2314 VSS nch l=0.04u w=0.4u
m4525 2334 2359 2315 VSS nch l=0.04u w=0.4u
m4526 70563 2206 VSS VSS nch l=0.04u w=0.8u
m4527 2336 2324 2316 VSS nch l=0.04u w=0.4u
m4528 2337 2267 2317 VSS nch l=0.04u w=0.4u
m4529 2338 2360 2318 VSS nch l=0.04u w=0.4u
m4530 70564 2210 VSS VSS nch l=0.04u w=0.8u
m4531 2340 FRAC[7] 2319 VSS nch l=0.04u w=0.4u
m4532 2341 2267 2320 VSS nch l=0.04u w=0.4u
m4533 2332 2295 2321 VSS nch l=0.04u w=0.4u
m4534 VSS 2252 VSS VSS nch l=0.26u w=0.8u
m4535 VSS 2255 VSS VSS nch l=0.26u w=0.8u
m4536 2349 2291 VSS VSS nch l=0.04u w=0.4u
m4537 2350 2292 VSS VSS nch l=0.04u w=0.4u
m4538 2351 2296 2322 VSS nch l=0.04u w=0.4u
m4539 2352 2297 2323 VSS nch l=0.04u w=0.4u
m4540 2353 2298 2324 VSS nch l=0.04u w=0.4u
m4541 2354 2299 2325 VSS nch l=0.04u w=0.4u
m4542 70566 2556 VSS VSS nch l=0.04u w=0.8u
m4543 70567 2557 VSS VSS nch l=0.04u w=0.8u
m4544 2357 2222 VSS VSS nch l=0.04u w=0.4u
m4545 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4546 70568 2289 VSS VSS nch l=0.04u w=0.24u
m4547 2326 2239 70560 VSS nch l=0.04u w=0.8u
m4548 2344 2308 2327 VSS nch l=0.04u w=0.4u
m4549 2328 2240 70561 VSS nch l=0.04u w=0.8u
m4550 2357 2309 2329 VSS nch l=0.04u w=0.4u
m4551 2330 2241 70562 VSS nch l=0.04u w=0.8u
m4552 FRAC[7] 2313 2331 VSS nch l=0.04u w=0.4u
m4553 2345 2314 2333 VSS nch l=0.04u w=0.4u
m4554 2359 2315 2334 VSS nch l=0.04u w=0.4u
m4555 2335 2242 70563 VSS nch l=0.04u w=0.8u
m4556 2324 2316 2336 VSS nch l=0.04u w=0.4u
m4557 2267 2317 2337 VSS nch l=0.04u w=0.4u
m4558 2360 2318 2338 VSS nch l=0.04u w=0.4u
m4559 2339 2243 70564 VSS nch l=0.04u w=0.8u
m4560 FRAC[7] 2319 2340 VSS nch l=0.04u w=0.4u
m4561 2267 2320 2341 VSS nch l=0.04u w=0.4u
m4562 2361 4328 VSS VSS nch l=0.04u w=0.4u
m4563 2362 4328 VSS VSS nch l=0.04u w=0.4u
m4564 2363 4328 VSS VSS nch l=0.04u w=0.4u
m4565 2364 4328 VSS VSS nch l=0.04u w=0.4u
m4566 2365 4328 VSS VSS nch l=0.04u w=0.4u
m4567 2366 4328 VSS VSS nch l=0.04u w=0.4u
m4568 70569 4328 2332 VSS nch l=0.04u w=0.12u
m4569 70573 4328 2351 VSS nch l=0.04u w=0.12u
m4570 70574 4328 2352 VSS nch l=0.04u w=0.12u
m4571 70575 4328 2353 VSS nch l=0.04u w=0.12u
m4572 70576 4328 2354 VSS nch l=0.04u w=0.12u
m4573 2355 3012 70566 VSS nch l=0.04u w=0.8u
m4574 2356 303 70567 VSS nch l=0.04u w=0.8u
m4575 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4576 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4577 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4578 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4579 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4580 2369 2454 70568 VSS nch l=0.04u w=0.24u
m4581 VSS 2252 VSS VSS nch l=0.26u w=0.8u
m4582 VSS 2255 VSS VSS nch l=0.26u w=0.8u
m4583 VSS 2381 70569 VSS nch l=0.04u w=0.12u
m4584 VSS 2349 2367 VSS nch l=0.04u w=0.4u
m4585 VSS 2350 2368 VSS nch l=0.04u w=0.4u
m4586 VSS 2392 70573 VSS nch l=0.04u w=0.12u
m4587 VSS 2393 70574 VSS nch l=0.04u w=0.12u
m4588 VSS 2394 70575 VSS nch l=0.04u w=0.12u
m4589 VSS 2395 70576 VSS nch l=0.04u w=0.12u
m4590 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4591 2188 2403 2369 VSS nch l=0.04u w=0.4u
m4592 70592 2302 2370 VSS nch l=0.04u w=0.8u
m4593 70593 2303 2371 VSS nch l=0.04u w=0.8u
m4594 2381 2332 VSS VSS nch l=0.04u w=0.4u
m4595 2375 2361 2373 VSS nch l=0.04u w=0.4u
m4596 2376 2362 2374 VSS nch l=0.04u w=0.4u
m4597 2377 2363 296 VSS nch l=0.04u w=0.4u
m4598 2378 2364 2310 VSS nch l=0.04u w=0.4u
m4599 2379 2365 2311 VSS nch l=0.04u w=0.4u
m4600 2380 2366 2312 VSS nch l=0.04u w=0.4u
m4601 710 2367 VSS VSS nch l=0.04u w=0.4u
m4602 1086 2368 VSS VSS nch l=0.04u w=0.4u
m4603 2392 2351 VSS VSS nch l=0.04u w=0.4u
m4604 2393 2352 VSS VSS nch l=0.04u w=0.4u
m4605 2394 2353 VSS VSS nch l=0.04u w=0.4u
m4606 2395 2354 VSS VSS nch l=0.04u w=0.4u
m4607 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4608 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4609 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4610 2396 2300 VSS VSS nch l=0.04u w=0.4u
m4611 2397 2301 VSS VSS nch l=0.04u w=0.4u
m4612 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4613 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4614 VSS 2252 VSS VSS nch l=0.26u w=0.8u
m4615 VSS 2255 VSS VSS nch l=0.26u w=0.8u
m4616 VSS 2143 70592 VSS nch l=0.04u w=0.8u
m4617 VSS 2147 70593 VSS nch l=0.04u w=0.8u
m4618 70595 4328 2375 VSS nch l=0.04u w=0.12u
m4619 70596 4328 2376 VSS nch l=0.04u w=0.12u
m4620 70597 4328 2377 VSS nch l=0.04u w=0.12u
m4621 2239 2405 2222 VSS nch l=0.04u w=0.4u
m4622 70598 2327 2382 VSS nch l=0.04u w=0.8u
m4623 2240 2406 139 VSS nch l=0.04u w=0.4u
m4624 70599 2329 2383 VSS nch l=0.04u w=0.8u
m4625 70600 4328 2378 VSS nch l=0.04u w=0.12u
m4626 70601 4328 2379 VSS nch l=0.04u w=0.12u
m4627 70602 4328 2380 VSS nch l=0.04u w=0.12u
m4628 2241 2407 FRAC[17] VSS nch l=0.04u w=0.4u
m4629 70603 2331 2384 VSS nch l=0.04u w=0.8u
m4630 70604 2333 2385 VSS nch l=0.04u w=0.8u
m4631 70605 2334 2386 VSS nch l=0.04u w=0.8u
m4632 2242 2408 1815 VSS nch l=0.04u w=0.4u
m4633 70606 2336 2387 VSS nch l=0.04u w=0.8u
m4634 70607 2337 2388 VSS nch l=0.04u w=0.8u
m4635 70608 2338 2389 VSS nch l=0.04u w=0.8u
m4636 2243 2409 FRAC[17] VSS nch l=0.04u w=0.4u
m4637 70609 2340 2390 VSS nch l=0.04u w=0.8u
m4638 70610 2341 2391 VSS nch l=0.04u w=0.8u
m4639 2398 155 VSS VSS nch l=0.04u w=0.4u
m4640 VSS 2300 2396 VSS nch l=0.04u w=0.4u
m4641 VSS 2301 2397 VSS nch l=0.04u w=0.4u
m4642 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4643 2400 2399 VSS VSS nch l=0.04u w=0.8u
m4644 2401 2402 VSS VSS nch l=0.04u w=0.8u
m4645 2403 2454 VSS VSS nch l=0.04u w=0.4u
m4646 VSS 2418 70595 VSS nch l=0.04u w=0.12u
m4647 VSS 2419 70596 VSS nch l=0.04u w=0.12u
m4648 VSS 2420 70597 VSS nch l=0.04u w=0.12u
m4649 2405 2222 2239 VSS nch l=0.04u w=0.4u
m4650 VSS 2159 70598 VSS nch l=0.04u w=0.8u
m4651 2406 139 2240 VSS nch l=0.04u w=0.4u
m4652 VSS 2161 70599 VSS nch l=0.04u w=0.8u
m4653 VSS 2422 70600 VSS nch l=0.04u w=0.12u
m4654 VSS 2423 70601 VSS nch l=0.04u w=0.12u
m4655 VSS 2424 70602 VSS nch l=0.04u w=0.12u
m4656 2407 FRAC[17] 2241 VSS nch l=0.04u w=0.4u
m4657 VSS 2163 70603 VSS nch l=0.04u w=0.8u
m4658 2404 4328 2381 VSS nch l=0.04u w=0.4u
m4659 VSS 2164 70604 VSS nch l=0.04u w=0.8u
m4660 VSS 2165 70605 VSS nch l=0.04u w=0.8u
m4661 2408 1815 2242 VSS nch l=0.04u w=0.4u
m4662 VSS 2167 70606 VSS nch l=0.04u w=0.8u
m4663 VSS 2168 70607 VSS nch l=0.04u w=0.8u
m4664 VSS 2169 70608 VSS nch l=0.04u w=0.8u
m4665 2409 FRAC[17] 2243 VSS nch l=0.04u w=0.4u
m4666 VSS 2171 70609 VSS nch l=0.04u w=0.8u
m4667 VSS 2172 70610 VSS nch l=0.04u w=0.8u
m4668 2410 4328 VSS VSS nch l=0.04u w=0.4u
m4669 2411 4328 VSS VSS nch l=0.04u w=0.4u
m4670 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4671 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4672 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4673 2412 4328 2392 VSS nch l=0.04u w=0.4u
m4674 2413 4328 2393 VSS nch l=0.04u w=0.4u
m4675 2414 4328 2394 VSS nch l=0.04u w=0.4u
m4676 2415 4328 2395 VSS nch l=0.04u w=0.4u
m4677 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4678 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4679 70612 2370 VSS VSS nch l=0.04u w=0.8u
m4680 2418 2375 VSS VSS nch l=0.04u w=0.4u
m4681 2419 2376 VSS VSS nch l=0.04u w=0.4u
m4682 2420 2377 VSS VSS nch l=0.04u w=0.4u
m4683 VSS 395 2405 VSS nch l=0.04u w=0.4u
m4684 70613 2371 VSS VSS nch l=0.04u w=0.8u
m4685 VSS 2225 2406 VSS nch l=0.04u w=0.4u
m4686 2422 2378 VSS VSS nch l=0.04u w=0.4u
m4687 2423 2379 VSS VSS nch l=0.04u w=0.4u
m4688 2424 2380 VSS VSS nch l=0.04u w=0.4u
m4689 VSS 2222 2407 VSS nch l=0.04u w=0.4u
m4690 70614 2295 2404 VSS nch l=0.04u w=0.12u
m4691 VSS 1941 2408 VSS nch l=0.04u w=0.4u
m4692 VSS 1942 2409 VSS nch l=0.04u w=0.4u
m4693 70617 155 VSS VSS nch l=0.04u w=0.8u
m4694 70618 2296 2412 VSS nch l=0.04u w=0.12u
m4695 70619 2297 2413 VSS nch l=0.04u w=0.12u
m4696 70620 2298 2414 VSS nch l=0.04u w=0.12u
m4697 70621 2299 2415 VSS nch l=0.04u w=0.12u
m4698 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4699 2426 2396 VSS VSS nch l=0.04u w=0.4u
m4700 2427 2397 VSS VSS nch l=0.04u w=0.4u
m4701 VSS 2454 2416 VSS nch l=0.04u w=0.4u
m4702 2417 2261 70612 VSS nch l=0.04u w=0.8u
m4703 2421 2262 70613 VSS nch l=0.04u w=0.8u
m4704 VSS 2453 70614 VSS nch l=0.04u w=0.12u
m4705 70623 2382 VSS VSS nch l=0.04u w=0.8u
m4706 70624 2383 VSS VSS nch l=0.04u w=0.8u
m4707 70625 2384 VSS VSS nch l=0.04u w=0.8u
m4708 70626 2385 VSS VSS nch l=0.04u w=0.8u
m4709 70627 2386 VSS VSS nch l=0.04u w=0.8u
m4710 70628 2387 VSS VSS nch l=0.04u w=0.8u
m4711 70629 2388 VSS VSS nch l=0.04u w=0.8u
m4712 70630 2389 VSS VSS nch l=0.04u w=0.8u
m4713 70631 2390 VSS VSS nch l=0.04u w=0.8u
m4714 70632 2391 VSS VSS nch l=0.04u w=0.8u
m4715 2425 FBDIV[7] 70617 VSS nch l=0.04u w=0.8u
m4716 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4717 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4718 VSS 2215 VSS VSS nch l=0.26u w=0.8u
m4719 2443 2410 2349 VSS nch l=0.04u w=0.4u
m4720 2444 2411 2350 VSS nch l=0.04u w=0.4u
m4721 VSS 2346 70618 VSS nch l=0.04u w=0.12u
m4722 VSS 2345 70619 VSS nch l=0.04u w=0.12u
m4723 VSS 2348 70620 VSS nch l=0.04u w=0.12u
m4724 VSS 2347 70621 VSS nch l=0.04u w=0.12u
m4725 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4726 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4727 VSS 2396 2426 VSS nch l=0.04u w=0.4u
m4728 VSS 2397 2427 VSS nch l=0.04u w=0.4u
m4729 2445 3454 VSS VSS nch l=0.04u w=0.4u
m4730 70634 2508 VSS VSS nch l=0.04u w=0.8u
m4731 2453 2404 VSS VSS nch l=0.04u w=0.4u
m4732 2447 4328 2418 VSS nch l=0.04u w=0.4u
m4733 2448 4328 2419 VSS nch l=0.04u w=0.4u
m4734 2449 4328 2420 VSS nch l=0.04u w=0.4u
m4735 70635 395 2428 VSS nch l=0.04u w=0.8u
m4736 2429 2272 70623 VSS nch l=0.04u w=0.8u
m4737 70636 2225 2430 VSS nch l=0.04u w=0.8u
m4738 2431 2273 70624 VSS nch l=0.04u w=0.8u
m4739 2450 4328 2422 VSS nch l=0.04u w=0.4u
m4740 2451 4328 2423 VSS nch l=0.04u w=0.4u
m4741 2452 4328 2424 VSS nch l=0.04u w=0.4u
m4742 70637 2222 2432 VSS nch l=0.04u w=0.8u
m4743 2433 2277 70625 VSS nch l=0.04u w=0.8u
m4744 2434 2278 70626 VSS nch l=0.04u w=0.8u
m4745 2435 2279 70627 VSS nch l=0.04u w=0.8u
m4746 70638 1941 2436 VSS nch l=0.04u w=0.8u
m4747 2437 2280 70628 VSS nch l=0.04u w=0.8u
m4748 2438 2281 70629 VSS nch l=0.04u w=0.8u
m4749 2439 2282 70630 VSS nch l=0.04u w=0.8u
m4750 70639 1942 2440 VSS nch l=0.04u w=0.8u
m4751 2441 2283 70631 VSS nch l=0.04u w=0.8u
m4752 2442 2284 70632 VSS nch l=0.04u w=0.8u
m4753 2455 2456 VSS VSS nch l=0.04u w=0.8u
m4754 70640 4328 2443 VSS nch l=0.04u w=0.12u
m4755 70641 4328 2444 VSS nch l=0.04u w=0.12u
m4756 VSS 2229 VSS VSS nch l=0.26u w=0.8u
m4757 2346 2412 VSS VSS nch l=0.04u w=0.4u
m4758 2345 2413 VSS VSS nch l=0.04u w=0.4u
m4759 2348 2414 VSS VSS nch l=0.04u w=0.4u
m4760 2347 2415 VSS VSS nch l=0.04u w=0.4u
m4761 2426 2396 VSS VSS nch l=0.04u w=0.4u
m4762 2427 2397 VSS VSS nch l=0.04u w=0.4u
m4763 2446 1918 70634 VSS nch l=0.04u w=0.8u
m4764 70643 2487 2454 VSS nch l=0.04u w=0.8u
m4765 2457 2302 VSS VSS nch l=0.04u w=0.4u
m4766 70644 2361 2447 VSS nch l=0.04u w=0.12u
m4767 70645 2362 2448 VSS nch l=0.04u w=0.12u
m4768 70646 2363 2449 VSS nch l=0.04u w=0.12u
m4769 VSS 2222 70635 VSS nch l=0.04u w=0.8u
m4770 2458 2303 VSS VSS nch l=0.04u w=0.4u
m4771 VSS 139 70636 VSS nch l=0.04u w=0.8u
m4772 70647 2364 2450 VSS nch l=0.04u w=0.12u
m4773 70648 2365 2451 VSS nch l=0.04u w=0.12u
m4774 70649 2366 2452 VSS nch l=0.04u w=0.12u
m4775 VSS FRAC[17] 70637 VSS nch l=0.04u w=0.8u
m4776 VSS 1815 70638 VSS nch l=0.04u w=0.8u
m4777 VSS FRAC[17] 70639 VSS nch l=0.04u w=0.8u
m4778 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4779 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4780 70651 2398 VSS VSS nch l=0.04u w=0.8u
m4781 VSS 2481 70640 VSS nch l=0.04u w=0.12u
m4782 VSS 2482 70641 VSS nch l=0.04u w=0.12u
m4783 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4784 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4785 2463 2462 VSS VSS nch l=0.04u w=0.8u
m4786 VSS 2396 2426 VSS nch l=0.04u w=0.4u
m4787 VSS 2397 2427 VSS nch l=0.04u w=0.4u
m4788 VSS 2648 70643 VSS nch l=0.04u w=0.8u
m4789 70654 2445 VSS VSS nch l=0.04u w=0.8u
m4790 2465 2143 2457 VSS nch l=0.04u w=0.4u
m4791 VSS 91 70644 VSS nch l=0.04u w=0.12u
m4792 VSS 2342 70645 VSS nch l=0.04u w=0.12u
m4793 VSS 125 70646 VSS nch l=0.04u w=0.12u
m4794 1041 2147 2458 VSS nch l=0.04u w=0.4u
m4795 VSS 2486 70647 VSS nch l=0.04u w=0.12u
m4796 VSS 2344 70648 VSS nch l=0.04u w=0.12u
m4797 VSS 129 70649 VSS nch l=0.04u w=0.12u
m4798 2467 2327 VSS VSS nch l=0.04u w=0.4u
m4799 2469 2329 VSS VSS nch l=0.04u w=0.4u
m4800 2471 2331 VSS VSS nch l=0.04u w=0.4u
m4801 2472 2333 VSS VSS nch l=0.04u w=0.4u
m4802 2473 2334 VSS VSS nch l=0.04u w=0.4u
m4803 2475 2336 VSS VSS nch l=0.04u w=0.4u
m4804 2476 2337 VSS VSS nch l=0.04u w=0.4u
m4805 2477 2338 VSS VSS nch l=0.04u w=0.4u
m4806 2479 2340 VSS VSS nch l=0.04u w=0.4u
m4807 2480 2341 VSS VSS nch l=0.04u w=0.4u
m4808 2459 2453 70651 VSS nch l=0.04u w=0.8u
m4809 2481 2443 VSS VSS nch l=0.04u w=0.4u
m4810 2482 2444 VSS VSS nch l=0.04u w=0.4u
m4811 VSS 2460 2460 VSS nch l=0.04u w=0.8u
m4812 2426 2396 VSS VSS nch l=0.04u w=0.4u
m4813 2427 2397 VSS VSS nch l=0.04u w=0.4u
m4814 2464 1918 70654 VSS nch l=0.04u w=0.8u
m4815 2485 1918 VSS VSS nch l=0.04u w=0.4u
m4816 2143 2457 2465 VSS nch l=0.04u w=0.4u
m4817 91 2447 VSS VSS nch l=0.04u w=0.4u
m4818 2342 2448 VSS VSS nch l=0.04u w=0.4u
m4819 VSS 2264 VSS VSS nch l=0.26u w=0.8u
m4820 125 2449 VSS VSS nch l=0.04u w=0.4u
m4821 2147 2458 1041 VSS nch l=0.04u w=0.4u
m4822 2486 2450 VSS VSS nch l=0.04u w=0.4u
m4823 2344 2451 VSS VSS nch l=0.04u w=0.4u
m4824 VSS 2266 VSS VSS nch l=0.26u w=0.8u
m4825 129 2452 VSS VSS nch l=0.04u w=0.4u
m4826 2374 2159 2467 VSS nch l=0.04u w=0.4u
m4827 2489 2161 2469 VSS nch l=0.04u w=0.4u
m4828 2343 2163 2471 VSS nch l=0.04u w=0.4u
m4829 2321 2164 2472 VSS nch l=0.04u w=0.4u
m4830 2323 2165 2473 VSS nch l=0.04u w=0.4u
m4831 2322 2167 2475 VSS nch l=0.04u w=0.4u
m4832 2359 2168 2476 VSS nch l=0.04u w=0.4u
m4833 2325 2169 2477 VSS nch l=0.04u w=0.4u
m4834 2324 2171 2479 VSS nch l=0.04u w=0.4u
m4835 2360 2172 2480 VSS nch l=0.04u w=0.4u
m4836 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4837 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4838 VSS 2484 2484 VSS nch l=0.04u w=0.8u
m4839 VSS 2396 2426 VSS nch l=0.04u w=0.4u
m4840 VSS 2397 2427 VSS nch l=0.04u w=0.4u
m4841 2491 2508 2485 VSS nch l=0.04u w=0.4u
m4842 2492 2493 VSS VSS nch l=0.04u w=0.8u
m4843 2494 2495 VSS VSS nch l=0.04u w=0.8u
m4844 VSS 2524 2487 VSS nch l=0.04u w=0.4u
m4845 2159 2467 2374 VSS nch l=0.04u w=0.4u
m4846 2161 2469 2489 VSS nch l=0.04u w=0.4u
m4847 2163 2471 2343 VSS nch l=0.04u w=0.4u
m4848 2164 2472 2321 VSS nch l=0.04u w=0.4u
m4849 2165 2473 2323 VSS nch l=0.04u w=0.4u
m4850 2167 2475 2322 VSS nch l=0.04u w=0.4u
m4851 2168 2476 2359 VSS nch l=0.04u w=0.4u
m4852 2169 2477 2325 VSS nch l=0.04u w=0.4u
m4853 2171 2479 2324 VSS nch l=0.04u w=0.4u
m4854 2172 2480 2360 VSS nch l=0.04u w=0.4u
m4855 2373 2511 2466 VSS nch l=0.04u w=0.4u
m4856 2488 2512 2468 VSS nch l=0.04u w=0.4u
m4857 2490 2513 2470 VSS nch l=0.04u w=0.4u
m4858 2153 2518 2474 VSS nch l=0.04u w=0.4u
m4859 2155 2523 2478 VSS nch l=0.04u w=0.4u
m4860 70671 2459 VSS VSS nch l=0.04u w=0.8u
m4861 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m4862 2504 4328 2481 VSS nch l=0.04u w=0.4u
m4863 2505 4328 2482 VSS nch l=0.04u w=0.4u
m4864 2426 2396 VSS VSS nch l=0.04u w=0.4u
m4865 2427 2397 VSS VSS nch l=0.04u w=0.4u
m4866 2508 2485 2491 VSS nch l=0.04u w=0.4u
m4867 70679 2416 VSS VSS nch l=0.04u w=0.12u
m4868 2509 2464 VSS VSS nch l=0.04u w=0.4u
m4869 2510 4328 VSS VSS nch l=0.04u w=0.4u
m4870 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4871 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4872 2511 2466 2373 VSS nch l=0.04u w=0.4u
m4873 2512 2468 2488 VSS nch l=0.04u w=0.4u
m4874 2513 2470 2490 VSS nch l=0.04u w=0.4u
m4875 2518 2474 2153 VSS nch l=0.04u w=0.4u
m4876 2523 2478 2155 VSS nch l=0.04u w=0.4u
m4877 2501 2425 70671 VSS nch l=0.04u w=0.8u
m4878 VSS 2503 2503 VSS nch l=0.04u w=0.8u
m4879 70682 2410 2504 VSS nch l=0.04u w=0.12u
m4880 70683 2411 2505 VSS nch l=0.04u w=0.12u
m4881 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m4882 VSS 2396 2426 VSS nch l=0.04u w=0.4u
m4883 VSS 2397 2427 VSS nch l=0.04u w=0.4u
m4884 VSS 2506 2506 VSS nch l=0.04u w=0.8u
m4885 2524 2615 70679 VSS nch l=0.04u w=0.12u
m4886 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m4887 2525 2417 VSS VSS nch l=0.04u w=0.4u
m4888 VSS 2496 2511 VSS nch l=0.04u w=0.4u
m4889 2526 2421 VSS VSS nch l=0.04u w=0.4u
m4890 VSS 2497 2512 VSS nch l=0.04u w=0.4u
m4891 VSS 2498 2513 VSS nch l=0.04u w=0.4u
m4892 VSS 2515 2515 VSS nch l=0.04u w=0.8u
m4893 VSS 2516 2516 VSS nch l=0.04u w=0.8u
m4894 VSS 2499 2518 VSS nch l=0.04u w=0.4u
m4895 VSS 2520 2520 VSS nch l=0.04u w=0.8u
m4896 VSS 2521 2521 VSS nch l=0.04u w=0.8u
m4897 VSS 2500 2523 VSS nch l=0.04u w=0.4u
m4898 VSS 2554 70682 VSS nch l=0.04u w=0.12u
m4899 VSS 2555 70683 VSS nch l=0.04u w=0.12u
m4900 VSS 2305 VSS VSS nch l=0.26u w=0.8u
m4901 VSS 2306 VSS VSS nch l=0.26u w=0.8u
m4902 2541 5232 2524 VSS nch l=0.04u w=0.4u
m4903 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m4904 2542 2510 LOCK VSS nch l=0.04u w=0.4u
m4905 2544 2429 VSS VSS nch l=0.04u w=0.4u
m4906 2545 2431 VSS VSS nch l=0.04u w=0.4u
m4907 2546 2433 VSS VSS nch l=0.04u w=0.4u
m4908 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m4909 2547 2434 VSS VSS nch l=0.04u w=0.4u
m4910 2548 2435 VSS VSS nch l=0.04u w=0.4u
m4911 2549 2437 VSS VSS nch l=0.04u w=0.4u
m4912 2550 2438 VSS VSS nch l=0.04u w=0.4u
m4913 2551 2439 VSS VSS nch l=0.04u w=0.4u
m4914 2552 2441 VSS VSS nch l=0.04u w=0.4u
m4915 2553 2442 VSS VSS nch l=0.04u w=0.4u
m4916 2554 2504 VSS VSS nch l=0.04u w=0.4u
m4917 2555 2505 VSS VSS nch l=0.04u w=0.4u
m4918 VSS 2527 2527 VSS nch l=0.04u w=0.8u
m4919 VSS 2530 2530 VSS nch l=0.04u w=0.8u
m4920 VSS 2531 2531 VSS nch l=0.04u w=0.8u
m4921 VSS 2534 2534 VSS nch l=0.04u w=0.8u
m4922 VSS 2535 2535 VSS nch l=0.04u w=0.8u
m4923 VSS 2538 2538 VSS nch l=0.04u w=0.8u
m4924 VSS 2539 2539 VSS nch l=0.04u w=0.8u
m4925 70704 2716 VSS VSS nch l=0.04u w=0.8u
m4926 70705 2716 VSS VSS nch l=0.04u w=0.8u
m4927 VSS 2507 VSS VSS nch l=0.26u w=0.8u
m4928 2558 2559 VSS VSS nch l=0.04u w=0.8u
m4929 2561 2560 VSS VSS nch l=0.04u w=0.8u
m4930 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m4931 VSS 2514 VSS VSS nch l=0.26u w=0.8u
m4932 VSS 2517 VSS VSS nch l=0.26u w=0.8u
m4933 VSS 2519 VSS VSS nch l=0.26u w=0.8u
m4934 VSS 2522 VSS VSS nch l=0.26u w=0.8u
m4935 70706 2491 2543 VSS nch l=0.04u w=0.8u
m4936 70707 4328 2542 VSS nch l=0.04u w=0.12u
m4937 70708 1464 VSS VSS nch l=0.04u w=0.8u
m4938 70709 2669 2198 VSS nch l=0.04u w=0.8u
m4939 70710 1465 VSS VSS nch l=0.04u w=0.8u
m4940 70711 2670 2200 VSS nch l=0.04u w=0.8u
m4941 70712 2671 2202 VSS nch l=0.04u w=0.8u
m4942 70713 2672 2206 VSS nch l=0.04u w=0.8u
m4943 70714 2673 2210 VSS nch l=0.04u w=0.8u
m4944 2556 2270 70704 VSS nch l=0.04u w=0.8u
m4945 2557 2271 70705 VSS nch l=0.04u w=0.8u
m4946 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m4947 70717 2594 2541 VSS nch l=0.04u w=0.8u
m4948 VSS 2630 70706 VSS nch l=0.04u w=0.8u
m4949 VSS 2580 70707 VSS nch l=0.04u w=0.12u
m4950 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m4951 70718 1755 70708 VSS nch l=0.04u w=0.8u
m4952 VSS 2584 70709 VSS nch l=0.04u w=0.8u
m4953 70719 1756 70710 VSS nch l=0.04u w=0.8u
m4954 VSS 2585 70711 VSS nch l=0.04u w=0.8u
m4955 VSS 2586 70712 VSS nch l=0.04u w=0.8u
m4956 VSS 2587 70713 VSS nch l=0.04u w=0.8u
m4957 VSS 2588 70714 VSS nch l=0.04u w=0.8u
m4958 70721 1488 VSS VSS nch l=0.04u w=0.8u
m4959 70722 1489 VSS VSS nch l=0.04u w=0.8u
m4960 70723 1490 VSS VSS nch l=0.04u w=0.8u
m4961 70724 1492 VSS VSS nch l=0.04u w=0.8u
m4962 70725 1493 VSS VSS nch l=0.04u w=0.8u
m4963 70726 1494 VSS VSS nch l=0.04u w=0.8u
m4964 70727 1495 VSS VSS nch l=0.04u w=0.8u
m4965 70728 1496 VSS VSS nch l=0.04u w=0.8u
m4966 70729 1497 VSS VSS nch l=0.04u w=0.8u
m4967 70730 1498 VSS VSS nch l=0.04u w=0.8u
m4968 2578 4328 VSS VSS nch l=0.04u w=0.4u
m4969 2579 4328 VSS VSS nch l=0.04u w=0.4u
m4970 VSS 2528 VSS VSS nch l=0.26u w=0.8u
m4971 VSS 2529 VSS VSS nch l=0.26u w=0.8u
m4972 VSS 2532 VSS VSS nch l=0.26u w=0.8u
m4973 VSS 2533 VSS VSS nch l=0.26u w=0.8u
m4974 VSS 2536 VSS VSS nch l=0.26u w=0.8u
m4975 VSS 2537 VSS VSS nch l=0.26u w=0.8u
m4976 VSS 2540 VSS VSS nch l=0.26u w=0.8u
m4977 VSS 2507 VSS VSS nch l=0.26u w=0.8u
m4978 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m4979 VSS 2514 VSS VSS nch l=0.26u w=0.8u
m4980 VSS 2517 VSS VSS nch l=0.26u w=0.8u
m4981 VSS 2519 VSS VSS nch l=0.26u w=0.8u
m4982 VSS 2522 VSS VSS nch l=0.26u w=0.8u
m4983 VSS 2564 2564 VSS nch l=0.04u w=0.8u
m4984 VSS 2567 2567 VSS nch l=0.04u w=0.8u
m4985 VSS 2648 70717 VSS nch l=0.04u w=0.8u
m4986 2580 2542 VSS VSS nch l=0.04u w=0.4u
m4987 2562 2038 70718 VSS nch l=0.04u w=0.8u
m4988 2563 2039 70719 VSS nch l=0.04u w=0.8u
m4989 70734 1774 70721 VSS nch l=0.04u w=0.8u
m4990 70735 1776 70722 VSS nch l=0.04u w=0.8u
m4991 70736 1778 70723 VSS nch l=0.04u w=0.8u
m4992 70737 1780 70724 VSS nch l=0.04u w=0.8u
m4993 70738 1781 70725 VSS nch l=0.04u w=0.8u
m4994 70739 1783 70726 VSS nch l=0.04u w=0.8u
m4995 70740 1784 70727 VSS nch l=0.04u w=0.8u
m4996 70741 1785 70728 VSS nch l=0.04u w=0.8u
m4997 70742 1787 70729 VSS nch l=0.04u w=0.8u
m4998 70743 1788 70730 VSS nch l=0.04u w=0.8u
m4999 2581 4353 VSS VSS nch l=0.04u w=0.4u
m5000 2582 11 VSS VSS nch l=0.04u w=0.4u
m5001 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m5002 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m5003 70746 2541 VSS VSS nch l=0.04u w=0.24u
m5004 70747 2543 VSS VSS nch l=0.04u w=0.8u
m5005 70749 2466 VSS VSS nch l=0.04u w=0.8u
m5006 2568 2056 70734 VSS nch l=0.04u w=0.8u
m5007 70750 2468 VSS VSS nch l=0.04u w=0.8u
m5008 2569 2058 70735 VSS nch l=0.04u w=0.8u
m5009 70751 2470 VSS VSS nch l=0.04u w=0.8u
m5010 2570 2060 70736 VSS nch l=0.04u w=0.8u
m5011 2571 2062 70737 VSS nch l=0.04u w=0.8u
m5012 2572 2063 70738 VSS nch l=0.04u w=0.8u
m5013 70752 2474 VSS VSS nch l=0.04u w=0.8u
m5014 2573 2065 70739 VSS nch l=0.04u w=0.8u
m5015 2574 2066 70740 VSS nch l=0.04u w=0.8u
m5016 2575 2067 70741 VSS nch l=0.04u w=0.8u
m5017 70753 2478 VSS VSS nch l=0.04u w=0.8u
m5018 2576 2069 70742 VSS nch l=0.04u w=0.8u
m5019 2577 2070 70743 VSS nch l=0.04u w=0.8u
m5020 VSS 2528 VSS VSS nch l=0.26u w=0.8u
m5021 VSS 2529 VSS VSS nch l=0.26u w=0.8u
m5022 VSS 2532 VSS VSS nch l=0.26u w=0.8u
m5023 VSS 2533 VSS VSS nch l=0.26u w=0.8u
m5024 VSS 2536 VSS VSS nch l=0.26u w=0.8u
m5025 VSS 2537 VSS VSS nch l=0.26u w=0.8u
m5026 VSS 2540 VSS VSS nch l=0.26u w=0.8u
m5027 2589 2578 2554 VSS nch l=0.04u w=0.4u
m5028 2590 2579 2555 VSS nch l=0.04u w=0.4u
m5029 VSS 2507 VSS VSS nch l=0.26u w=0.8u
m5030 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m5031 VSS 2514 VSS VSS nch l=0.26u w=0.8u
m5032 VSS 2517 VSS VSS nch l=0.26u w=0.8u
m5033 VSS 2519 VSS VSS nch l=0.26u w=0.8u
m5034 VSS 2522 VSS VSS nch l=0.26u w=0.8u
m5035 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5036 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5037 2594 5232 70746 VSS nch l=0.04u w=0.24u
m5038 2583 2446 70747 VSS nch l=0.04u w=0.8u
m5039 2593 4328 2580 VSS nch l=0.04u w=0.4u
m5040 2595 2562 VSS VSS nch l=0.04u w=0.4u
m5041 2584 2496 70749 VSS nch l=0.04u w=0.8u
m5042 2596 2563 VSS VSS nch l=0.04u w=0.4u
m5043 2585 2497 70750 VSS nch l=0.04u w=0.8u
m5044 2586 2498 70751 VSS nch l=0.04u w=0.8u
m5045 2587 2499 70752 VSS nch l=0.04u w=0.8u
m5046 2588 2500 70753 VSS nch l=0.04u w=0.8u
m5047 70757 4328 2589 VSS nch l=0.04u w=0.12u
m5048 70758 4328 2590 VSS nch l=0.04u w=0.12u
m5049 VSS 2592 2592 VSS nch l=0.04u w=0.8u
m5050 2597 2581 2355 VSS nch l=0.04u w=0.4u
m5051 2598 2582 2356 VSS nch l=0.04u w=0.4u
m5052 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m5053 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m5054 2454 2615 2594 VSS nch l=0.04u w=0.4u
m5055 70761 2510 2593 VSS nch l=0.04u w=0.12u
m5056 VSS 2528 VSS VSS nch l=0.26u w=0.8u
m5057 VSS 2529 VSS VSS nch l=0.26u w=0.8u
m5058 VSS 2532 VSS VSS nch l=0.26u w=0.8u
m5059 VSS 2533 VSS VSS nch l=0.26u w=0.8u
m5060 VSS 2536 VSS VSS nch l=0.26u w=0.8u
m5061 VSS 2537 VSS VSS nch l=0.26u w=0.8u
m5062 VSS 2540 VSS VSS nch l=0.26u w=0.8u
m5063 2599 2568 VSS VSS nch l=0.04u w=0.4u
m5064 2600 2569 VSS VSS nch l=0.04u w=0.4u
m5065 2602 2570 VSS VSS nch l=0.04u w=0.4u
m5066 2603 2571 VSS VSS nch l=0.04u w=0.4u
m5067 2604 2572 VSS VSS nch l=0.04u w=0.4u
m5068 2605 2573 VSS VSS nch l=0.04u w=0.4u
m5069 2606 2574 VSS VSS nch l=0.04u w=0.4u
m5070 2607 2575 VSS VSS nch l=0.04u w=0.4u
m5071 2608 2576 VSS VSS nch l=0.04u w=0.4u
m5072 2609 2577 VSS VSS nch l=0.04u w=0.4u
m5073 VSS 2613 70757 VSS nch l=0.04u w=0.12u
m5074 VSS 2614 70758 VSS nch l=0.04u w=0.12u
m5075 VSS 2507 VSS VSS nch l=0.26u w=0.8u
m5076 70768 4353 2597 VSS nch l=0.04u w=0.12u
m5077 70769 11 2598 VSS nch l=0.04u w=0.12u
m5078 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m5079 VSS 2514 VSS VSS nch l=0.26u w=0.8u
m5080 VSS 2517 VSS VSS nch l=0.26u w=0.8u
m5081 VSS 2519 VSS VSS nch l=0.26u w=0.8u
m5082 VSS 2522 VSS VSS nch l=0.26u w=0.8u
m5083 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5084 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5085 VSS 2616 70761 VSS nch l=0.04u w=0.12u
m5086 2610 2491 VSS VSS nch l=0.04u w=0.4u
m5087 70770 2595 VSS VSS nch l=0.04u w=0.8u
m5088 70771 2596 VSS VSS nch l=0.04u w=0.8u
m5089 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5090 2613 2589 VSS VSS nch l=0.04u w=0.4u
m5091 2614 2590 VSS VSS nch l=0.04u w=0.4u
m5092 VSS 2628 70768 VSS nch l=0.04u w=0.12u
m5093 VSS 2629 70769 VSS nch l=0.04u w=0.12u
m5094 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m5095 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m5096 2615 5232 VSS VSS nch l=0.04u w=0.4u
m5097 VSS 2528 VSS VSS nch l=0.26u w=0.8u
m5098 VSS 2529 VSS VSS nch l=0.26u w=0.8u
m5099 VSS 2532 VSS VSS nch l=0.26u w=0.8u
m5100 VSS 2533 VSS VSS nch l=0.26u w=0.8u
m5101 VSS 2536 VSS VSS nch l=0.26u w=0.8u
m5102 VSS 2537 VSS VSS nch l=0.26u w=0.8u
m5103 VSS 2540 VSS VSS nch l=0.26u w=0.8u
m5104 2616 2593 VSS VSS nch l=0.04u w=0.4u
m5105 2617 2630 2610 VSS nch l=0.04u w=0.4u
m5106 70773 2302 70770 VSS nch l=0.04u w=0.8u
m5107 70774 2303 70771 VSS nch l=0.04u w=0.8u
m5108 VSS 2507 VSS VSS nch l=0.26u w=0.8u
m5109 2496 2633 2486 VSS nch l=0.04u w=0.4u
m5110 70775 2599 VSS VSS nch l=0.04u w=0.8u
m5111 2497 2634 2097 VSS nch l=0.04u w=0.4u
m5112 70776 2600 VSS VSS nch l=0.04u w=0.8u
m5113 2498 2635 FRAC[16] VSS nch l=0.04u w=0.4u
m5114 70777 2602 VSS VSS nch l=0.04u w=0.8u
m5115 70778 2603 VSS VSS nch l=0.04u w=0.8u
m5116 70779 2604 VSS VSS nch l=0.04u w=0.8u
m5117 2499 2638 2155 VSS nch l=0.04u w=0.4u
m5118 70780 2605 VSS VSS nch l=0.04u w=0.8u
m5119 70781 2606 VSS VSS nch l=0.04u w=0.8u
m5120 70782 2607 VSS VSS nch l=0.04u w=0.8u
m5121 2500 2639 FRAC[16] VSS nch l=0.04u w=0.4u
m5122 70783 2608 VSS VSS nch l=0.04u w=0.8u
m5123 70784 2609 VSS VSS nch l=0.04u w=0.8u
m5124 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m5125 VSS 2514 VSS VSS nch l=0.26u w=0.8u
m5126 VSS 2517 VSS VSS nch l=0.26u w=0.8u
m5127 VSS 2519 VSS VSS nch l=0.26u w=0.8u
m5128 VSS 2522 VSS VSS nch l=0.26u w=0.8u
m5129 2628 2597 VSS VSS nch l=0.04u w=0.4u
m5130 2629 2598 VSS VSS nch l=0.04u w=0.4u
m5131 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5132 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5133 2630 2610 2617 VSS nch l=0.04u w=0.4u
m5134 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5135 2611 1370 70773 VSS nch l=0.04u w=0.8u
m5136 2612 1371 70774 VSS nch l=0.04u w=0.8u
m5137 2631 2632 VSS VSS nch l=0.04u w=0.8u
m5138 2633 2486 2496 VSS nch l=0.04u w=0.4u
m5139 70785 2327 70775 VSS nch l=0.04u w=0.8u
m5140 2634 2097 2497 VSS nch l=0.04u w=0.4u
m5141 70786 2329 70776 VSS nch l=0.04u w=0.8u
m5142 2635 FRAC[16] 2498 VSS nch l=0.04u w=0.4u
m5143 70787 2331 70777 VSS nch l=0.04u w=0.8u
m5144 70788 2333 70778 VSS nch l=0.04u w=0.8u
m5145 70789 2334 70779 VSS nch l=0.04u w=0.8u
m5146 2638 2155 2499 VSS nch l=0.04u w=0.4u
m5147 70790 2336 70780 VSS nch l=0.04u w=0.8u
m5148 70791 2337 70781 VSS nch l=0.04u w=0.8u
m5149 70792 2338 70782 VSS nch l=0.04u w=0.8u
m5150 2639 FRAC[16] 2500 VSS nch l=0.04u w=0.4u
m5151 70793 2340 70783 VSS nch l=0.04u w=0.8u
m5152 70794 2341 70784 VSS nch l=0.04u w=0.8u
m5153 2636 4328 2613 VSS nch l=0.04u w=0.4u
m5154 2637 4328 2614 VSS nch l=0.04u w=0.4u
m5155 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m5156 2641 2640 VSS VSS nch l=0.04u w=0.8u
m5157 2642 2643 VSS VSS nch l=0.04u w=0.8u
m5158 2645 2644 VSS VSS nch l=0.04u w=0.8u
m5159 2646 2647 VSS VSS nch l=0.04u w=0.8u
m5160 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m5161 VSS 2528 VSS VSS nch l=0.26u w=0.8u
m5162 VSS 2529 VSS VSS nch l=0.26u w=0.8u
m5163 VSS 2532 VSS VSS nch l=0.26u w=0.8u
m5164 VSS 2533 VSS VSS nch l=0.26u w=0.8u
m5165 VSS 2536 VSS VSS nch l=0.26u w=0.8u
m5166 VSS 2537 VSS VSS nch l=0.26u w=0.8u
m5167 VSS 2540 VSS VSS nch l=0.26u w=0.8u
m5168 2648 2759 VSS VSS nch l=0.04u w=0.4u
m5169 2649 2649 VSS VSS nch l=0.04u w=0.8u
m5170 VSS 91 2633 VSS nch l=0.04u w=0.4u
m5171 2618 1380 70785 VSS nch l=0.04u w=0.8u
m5172 VSS 2490 2634 VSS nch l=0.04u w=0.4u
m5173 2619 1382 70786 VSS nch l=0.04u w=0.8u
m5174 VSS 2486 2635 VSS nch l=0.04u w=0.4u
m5175 2620 1384 70787 VSS nch l=0.04u w=0.8u
m5176 2621 1385 70788 VSS nch l=0.04u w=0.8u
m5177 2622 1386 70789 VSS nch l=0.04u w=0.8u
m5178 VSS 2287 2638 VSS nch l=0.04u w=0.4u
m5179 2623 1387 70790 VSS nch l=0.04u w=0.8u
m5180 2624 1388 70791 VSS nch l=0.04u w=0.8u
m5181 2625 1389 70792 VSS nch l=0.04u w=0.8u
m5182 VSS 2288 2639 VSS nch l=0.04u w=0.4u
m5183 2626 1390 70793 VSS nch l=0.04u w=0.8u
m5184 2627 1391 70794 VSS nch l=0.04u w=0.8u
m5185 70795 2578 2636 VSS nch l=0.04u w=0.12u
m5186 70796 2579 2637 VSS nch l=0.04u w=0.12u
m5187 VSS 2461 VSS VSS nch l=0.26u w=0.8u
m5188 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5189 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5190 2650 4353 2628 VSS nch l=0.04u w=0.4u
m5191 2651 11 2629 VSS nch l=0.04u w=0.4u
m5192 2652 2653 VSS VSS nch l=0.04u w=0.8u
m5193 2655 2654 VSS VSS nch l=0.04u w=0.8u
m5194 2656 2657 VSS VSS nch l=0.04u w=0.8u
m5195 2659 2658 VSS VSS nch l=0.04u w=0.8u
m5196 2660 2661 VSS VSS nch l=0.04u w=0.8u
m5197 2663 2662 VSS VSS nch l=0.04u w=0.8u
m5198 2664 2665 VSS VSS nch l=0.04u w=0.8u
m5199 VSS 2759 2648 VSS nch l=0.04u w=0.4u
m5200 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5201 2666 2445 VSS VSS nch l=0.04u w=0.4u
m5202 70799 2525 VSS VSS nch l=0.04u w=0.8u
m5203 70800 2526 VSS VSS nch l=0.04u w=0.8u
m5204 VSS 2681 70795 VSS nch l=0.04u w=0.12u
m5205 VSS 2682 70796 VSS nch l=0.04u w=0.12u
m5206 2674 2675 VSS VSS nch l=0.04u w=0.8u
m5207 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m5208 VSS 2483 VSS VSS nch l=0.26u w=0.8u
m5209 70801 2581 2650 VSS nch l=0.04u w=0.12u
m5210 70802 2582 2651 VSS nch l=0.04u w=0.12u
m5211 315 2676 VSS VSS nch l=0.04u w=0.8u
m5212 VSS 2617 2666 VSS nch l=0.04u w=0.4u
m5213 70803 2508 VSS VSS nch l=0.04u w=0.8u
m5214 2667 2611 70799 VSS nch l=0.04u w=0.8u
m5215 2668 2612 70800 VSS nch l=0.04u w=0.8u
m5216 70804 91 2669 VSS nch l=0.04u w=0.8u
m5217 70805 2544 VSS VSS nch l=0.04u w=0.8u
m5218 70806 2490 2670 VSS nch l=0.04u w=0.8u
m5219 70807 2545 VSS VSS nch l=0.04u w=0.8u
m5220 70808 2486 2671 VSS nch l=0.04u w=0.8u
m5221 70809 2546 VSS VSS nch l=0.04u w=0.8u
m5222 2681 2636 VSS VSS nch l=0.04u w=0.4u
m5223 2682 2637 VSS VSS nch l=0.04u w=0.4u
m5224 70810 2547 VSS VSS nch l=0.04u w=0.8u
m5225 70811 2548 VSS VSS nch l=0.04u w=0.8u
m5226 70812 2287 2672 VSS nch l=0.04u w=0.8u
m5227 70813 2549 VSS VSS nch l=0.04u w=0.8u
m5228 70814 2550 VSS VSS nch l=0.04u w=0.8u
m5229 70815 2551 VSS VSS nch l=0.04u w=0.8u
m5230 70816 2288 2673 VSS nch l=0.04u w=0.8u
m5231 70817 2552 VSS VSS nch l=0.04u w=0.8u
m5232 70818 2553 VSS VSS nch l=0.04u w=0.8u
m5233 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5234 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5235 2693 2692 VSS VSS nch l=0.04u w=0.8u
m5236 VSS 2696 70801 VSS nch l=0.04u w=0.12u
m5237 VSS 2697 70802 VSS nch l=0.04u w=0.12u
m5238 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5239 2677 2197 70803 VSS nch l=0.04u w=0.8u
m5240 VSS 2486 70804 VSS nch l=0.04u w=0.8u
m5241 2678 2618 70805 VSS nch l=0.04u w=0.8u
m5242 VSS 2502 VSS VSS nch l=0.26u w=0.8u
m5243 VSS 2097 70806 VSS nch l=0.04u w=0.8u
m5244 2679 2619 70807 VSS nch l=0.04u w=0.8u
m5245 VSS FRAC[16] 70808 VSS nch l=0.04u w=0.8u
m5246 2680 2620 70809 VSS nch l=0.04u w=0.8u
m5247 2683 2621 70810 VSS nch l=0.04u w=0.8u
m5248 2684 2622 70811 VSS nch l=0.04u w=0.8u
m5249 VSS 2155 70812 VSS nch l=0.04u w=0.8u
m5250 2685 2623 70813 VSS nch l=0.04u w=0.8u
m5251 2686 2624 70814 VSS nch l=0.04u w=0.8u
m5252 2687 2625 70815 VSS nch l=0.04u w=0.8u
m5253 VSS FRAC[16] 70816 VSS nch l=0.04u w=0.8u
m5254 2688 2626 70817 VSS nch l=0.04u w=0.8u
m5255 2689 2627 70818 VSS nch l=0.04u w=0.8u
m5256 VSS 2690 2690 VSS nch l=0.04u w=0.8u
m5257 2696 2650 VSS VSS nch l=0.04u w=0.4u
m5258 2697 2651 VSS VSS nch l=0.04u w=0.4u
m5259 70834 2445 VSS VSS nch l=0.04u w=0.8u
m5260 70835 110 VSS VSS nch l=0.04u w=0.8u
m5261 2702 2702 VSS VSS nch l=0.04u w=0.8u
m5262 2704 2703 VSS VSS nch l=0.04u w=0.8u
m5263 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5264 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5265 2713 4328 VSS VSS nch l=0.04u w=0.4u
m5266 2714 4328 VSS VSS nch l=0.04u w=0.4u
m5267 VSS 2695 2695 VSS nch l=0.04u w=0.8u
m5268 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5269 VSS 2698 2698 VSS nch l=0.04u w=0.8u
m5270 2700 2197 70834 VSS nch l=0.04u w=0.8u
m5271 2717 2197 VSS VSS nch l=0.04u w=0.4u
m5272 2701 125 70835 VSS nch l=0.04u w=0.8u
m5273 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5274 VSS 2705 2705 VSS nch l=0.04u w=0.8u
m5275 VSS 2708 2708 VSS nch l=0.04u w=0.8u
m5276 70838 2753 2466 VSS nch l=0.04u w=0.8u
m5277 70839 2795 VSS VSS nch l=0.04u w=0.8u
m5278 70840 2754 2468 VSS nch l=0.04u w=0.8u
m5279 70841 1853 VSS VSS nch l=0.04u w=0.8u
m5280 70842 2616 VSS VSS nch l=0.04u w=0.8u
m5281 70843 2616 VSS VSS nch l=0.04u w=0.8u
m5282 VSS 2709 2709 VSS nch l=0.04u w=0.8u
m5283 VSS 2712 2712 VSS nch l=0.04u w=0.8u
m5284 70844 2755 2470 VSS nch l=0.04u w=0.8u
m5285 70845 FRAC[8] VSS VSS nch l=0.04u w=0.8u
m5286 VSS 2774 2715 VSS nch l=0.04u w=0.4u
m5287 70846 2796 VSS VSS nch l=0.04u w=0.8u
m5288 2728 4328 VSS VSS nch l=0.04u w=0.4u
m5289 2729 4328 VSS VSS nch l=0.04u w=0.4u
m5290 70847 2804 VSS VSS nch l=0.04u w=0.8u
m5291 70848 2757 2474 VSS nch l=0.04u w=0.8u
m5292 70849 2805 VSS VSS nch l=0.04u w=0.8u
m5293 70850 2715 VSS VSS nch l=0.04u w=0.8u
m5294 2733 4328 VSS VSS nch l=0.04u w=0.4u
m5295 2734 4328 VSS VSS nch l=0.04u w=0.4u
m5296 70851 2808 VSS VSS nch l=0.04u w=0.8u
m5297 70852 2758 2478 VSS nch l=0.04u w=0.8u
m5298 70853 FRAC[8] VSS VSS nch l=0.04u w=0.8u
m5299 70854 2715 VSS VSS nch l=0.04u w=0.8u
m5300 2738 PD VSS VSS nch l=0.04u w=0.4u
m5301 VSS 2746 2716 VSS nch l=0.04u w=0.4u
m5302 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5303 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5304 2739 2508 2717 VSS nch l=0.04u w=0.4u
m5305 VSS 2889 70838 VSS nch l=0.04u w=0.8u
m5306 2718 2793 70839 VSS nch l=0.04u w=0.8u
m5307 VSS 2719 2719 VSS nch l=0.04u w=0.8u
m5308 VSS 2722 2722 VSS nch l=0.04u w=0.8u
m5309 VSS 2890 70840 VSS nch l=0.04u w=0.8u
m5310 2723 2794 70841 VSS nch l=0.04u w=0.8u
m5311 2724 2928 70842 VSS nch l=0.04u w=0.8u
m5312 2725 2929 70843 VSS nch l=0.04u w=0.8u
m5313 VSS 2891 70844 VSS nch l=0.04u w=0.8u
m5314 2726 2795 70845 VSS nch l=0.04u w=0.8u
m5315 2727 131 70846 VSS nch l=0.04u w=0.8u
m5316 2730 2796 70847 VSS nch l=0.04u w=0.8u
m5317 VSS 2892 70848 VSS nch l=0.04u w=0.8u
m5318 2731 2797 70849 VSS nch l=0.04u w=0.8u
m5319 2732 2798 70850 VSS nch l=0.04u w=0.8u
m5320 2735 2799 70851 VSS nch l=0.04u w=0.8u
m5321 VSS 2893 70852 VSS nch l=0.04u w=0.8u
m5322 2736 2800 70853 VSS nch l=0.04u w=0.8u
m5323 2737 FBDIV[8] 70854 VSS nch l=0.04u w=0.8u
m5324 2740 2713 2681 VSS nch l=0.04u w=0.4u
m5325 2741 2714 2682 VSS nch l=0.04u w=0.4u
m5326 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5327 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5328 VSS 2699 VSS VSS nch l=0.26u w=0.8u
m5329 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5330 2508 2717 2739 VSS nch l=0.04u w=0.4u
m5331 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5332 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5333 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5334 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5335 2747 2700 VSS VSS nch l=0.04u w=0.4u
m5336 2748 125 VSS VSS nch l=0.04u w=0.4u
m5337 70859 4328 2740 VSS nch l=0.04u w=0.12u
m5338 70860 4328 2741 VSS nch l=0.04u w=0.12u
m5339 2756 4328 VSS VSS nch l=0.04u w=0.4u
m5340 2749 2728 2742 VSS nch l=0.04u w=0.4u
m5341 2750 2729 2743 VSS nch l=0.04u w=0.4u
m5342 2751 2733 2744 VSS nch l=0.04u w=0.4u
m5343 2752 2734 2745 VSS nch l=0.04u w=0.4u
m5344 70861 2738 VSS VSS nch l=0.04u w=0.8u
m5345 2760 5232 2746 VSS nch l=0.04u w=0.62u
m5346 VSS 2565 VSS VSS nch l=0.26u w=0.8u
m5347 VSS 2566 VSS VSS nch l=0.26u w=0.8u
m5348 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5349 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5350 2761 110 2748 VSS nch l=0.04u w=0.4u
m5351 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5352 70862 3737 2753 VSS nch l=0.04u w=0.8u
m5353 2762 2793 VSS VSS nch l=0.04u w=0.4u
m5354 70863 3739 2754 VSS nch l=0.04u w=0.8u
m5355 2763 2794 VSS VSS nch l=0.04u w=0.4u
m5356 2764 2724 VSS VSS nch l=0.04u w=0.4u
m5357 2765 2725 VSS VSS nch l=0.04u w=0.4u
m5358 70864 3741 2755 VSS nch l=0.04u w=0.8u
m5359 2766 2795 VSS VSS nch l=0.04u w=0.4u
m5360 VSS 2783 70859 VSS nch l=0.04u w=0.12u
m5361 VSS 2784 70860 VSS nch l=0.04u w=0.12u
m5362 2767 131 VSS VSS nch l=0.04u w=0.4u
m5363 70865 4328 2749 VSS nch l=0.04u w=0.12u
m5364 70866 4328 2750 VSS nch l=0.04u w=0.12u
m5365 2768 2796 VSS VSS nch l=0.04u w=0.4u
m5366 70867 3745 2757 VSS nch l=0.04u w=0.8u
m5367 2769 2797 VSS VSS nch l=0.04u w=0.4u
m5368 2770 2798 VSS VSS nch l=0.04u w=0.4u
m5369 70868 4328 2751 VSS nch l=0.04u w=0.12u
m5370 70869 4328 2752 VSS nch l=0.04u w=0.12u
m5371 2771 2799 VSS VSS nch l=0.04u w=0.4u
m5372 70870 3749 2758 VSS nch l=0.04u w=0.8u
m5373 2772 2800 VSS VSS nch l=0.04u w=0.4u
m5374 2773 FBDIV[8] VSS VSS nch l=0.04u w=0.4u
m5375 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5376 70872 2696 70861 VSS nch l=0.04u w=0.8u
m5377 VSS 2738 2760 VSS nch l=0.04u w=0.8u
m5378 VSS 2699 VSS VSS nch l=0.26u w=0.8u
m5379 2775 2776 VSS VSS nch l=0.04u w=0.8u
m5380 2778 2777 VSS VSS nch l=0.04u w=0.8u
m5381 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5382 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5383 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5384 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5385 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5386 110 2748 2761 VSS nch l=0.04u w=0.4u
m5387 70873 2947 70862 VSS nch l=0.04u w=0.8u
m5388 2780 2795 2762 VSS nch l=0.04u w=0.4u
m5389 70874 2948 70863 VSS nch l=0.04u w=0.8u
m5390 2781 1853 2763 VSS nch l=0.04u w=0.4u
m5391 70875 2949 70864 VSS nch l=0.04u w=0.8u
m5392 2782 FRAC[8] 2766 VSS nch l=0.04u w=0.4u
m5393 2783 2740 VSS VSS nch l=0.04u w=0.4u
m5394 2784 2741 VSS VSS nch l=0.04u w=0.4u
m5395 2786 2796 2767 VSS nch l=0.04u w=0.4u
m5396 VSS 2802 70865 VSS nch l=0.04u w=0.12u
m5397 VSS 2803 70866 VSS nch l=0.04u w=0.12u
m5398 2787 2804 2768 VSS nch l=0.04u w=0.4u
m5399 70876 2950 70867 VSS nch l=0.04u w=0.8u
m5400 2788 2805 2769 VSS nch l=0.04u w=0.4u
m5401 2789 2715 2770 VSS nch l=0.04u w=0.4u
m5402 VSS 2806 70868 VSS nch l=0.04u w=0.12u
m5403 VSS 2807 70869 VSS nch l=0.04u w=0.12u
m5404 2790 2808 2771 VSS nch l=0.04u w=0.4u
m5405 70877 2951 70870 VSS nch l=0.04u w=0.8u
m5406 2791 FRAC[8] 2772 VSS nch l=0.04u w=0.4u
m5407 2792 2715 2773 VSS nch l=0.04u w=0.4u
m5408 2785 2756 2774 VSS nch l=0.04u w=0.4u
m5409 2759 2697 70872 VSS nch l=0.04u w=0.8u
m5410 2760 2738 VSS VSS nch l=0.04u w=0.8u
m5411 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5412 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5413 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5414 70878 2739 2779 VSS nch l=0.04u w=0.8u
m5415 VSS 2816 70873 VSS nch l=0.04u w=0.8u
m5416 2795 2762 2780 VSS nch l=0.04u w=0.4u
m5417 VSS 2817 70874 VSS nch l=0.04u w=0.8u
m5418 1853 2763 2781 VSS nch l=0.04u w=0.4u
m5419 VSS 2818 70875 VSS nch l=0.04u w=0.8u
m5420 FRAC[8] 2766 2782 VSS nch l=0.04u w=0.4u
m5421 2796 2767 2786 VSS nch l=0.04u w=0.4u
m5422 2802 2749 VSS VSS nch l=0.04u w=0.4u
m5423 2803 2750 VSS VSS nch l=0.04u w=0.4u
m5424 2804 2768 2787 VSS nch l=0.04u w=0.4u
m5425 VSS 2819 70876 VSS nch l=0.04u w=0.8u
m5426 2805 2769 2788 VSS nch l=0.04u w=0.4u
m5427 2715 2770 2789 VSS nch l=0.04u w=0.4u
m5428 2806 2751 VSS VSS nch l=0.04u w=0.4u
m5429 2807 2752 VSS VSS nch l=0.04u w=0.4u
m5430 2808 2771 2790 VSS nch l=0.04u w=0.4u
m5431 VSS 2820 70877 VSS nch l=0.04u w=0.8u
m5432 FRAC[8] 2772 2791 VSS nch l=0.04u w=0.4u
m5433 2715 2773 2792 VSS nch l=0.04u w=0.4u
m5434 2809 4328 VSS VSS nch l=0.04u w=0.4u
m5435 2810 4328 VSS VSS nch l=0.04u w=0.4u
m5436 2811 4328 VSS VSS nch l=0.04u w=0.4u
m5437 2812 4328 VSS VSS nch l=0.04u w=0.4u
m5438 70881 4328 2785 VSS nch l=0.04u w=0.12u
m5439 VSS 2591 VSS VSS nch l=0.26u w=0.8u
m5440 VSS 2699 VSS VSS nch l=0.26u w=0.8u
m5441 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5442 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5443 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5444 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5445 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5446 VSS 2583 70878 VSS nch l=0.04u w=0.8u
m5447 2813 4328 2783 VSS nch l=0.04u w=0.4u
m5448 2814 4328 2784 VSS nch l=0.04u w=0.4u
m5449 VSS 2833 70881 VSS nch l=0.04u w=0.12u
m5450 2822 2821 VSS VSS nch l=0.04u w=0.8u
m5451 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5452 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5453 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5454 70895 2761 2815 VSS nch l=0.04u w=0.8u
m5455 VSS 2845 2816 VSS nch l=0.04u w=0.4u
m5456 VSS 2846 2817 VSS nch l=0.04u w=0.4u
m5457 VSS 2847 2818 VSS nch l=0.04u w=0.4u
m5458 70896 2713 2813 VSS nch l=0.04u w=0.12u
m5459 70897 2714 2814 VSS nch l=0.04u w=0.12u
m5460 2833 2785 VSS VSS nch l=0.04u w=0.4u
m5461 2825 4328 2802 VSS nch l=0.04u w=0.4u
m5462 2826 4328 2803 VSS nch l=0.04u w=0.4u
m5463 VSS 2848 2819 VSS nch l=0.04u w=0.4u
m5464 2827 4328 2806 VSS nch l=0.04u w=0.4u
m5465 2828 4328 2807 VSS nch l=0.04u w=0.4u
m5466 VSS 2849 2820 VSS nch l=0.04u w=0.4u
m5467 2829 2809 2823 VSS nch l=0.04u w=0.4u
m5468 2830 2810 2824 VSS nch l=0.04u w=0.4u
m5469 2831 2811 2764 VSS nch l=0.04u w=0.4u
m5470 2832 2812 2765 VSS nch l=0.04u w=0.4u
m5471 VSS 2699 VSS VSS nch l=0.26u w=0.8u
m5472 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5473 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5474 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5475 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5476 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5477 70902 2779 VSS VSS nch l=0.04u w=0.8u
m5478 VSS 2667 70895 VSS nch l=0.04u w=0.8u
m5479 VSS 2851 70896 VSS nch l=0.04u w=0.12u
m5480 VSS 2852 70897 VSS nch l=0.04u w=0.12u
m5481 70903 2728 2825 VSS nch l=0.04u w=0.12u
m5482 70904 2729 2826 VSS nch l=0.04u w=0.12u
m5483 70905 2733 2827 VSS nch l=0.04u w=0.12u
m5484 70906 2734 2828 VSS nch l=0.04u w=0.12u
m5485 70908 4328 2829 VSS nch l=0.04u w=0.12u
m5486 70909 4328 2830 VSS nch l=0.04u w=0.12u
m5487 70910 2780 2834 VSS nch l=0.04u w=0.8u
m5488 70911 2781 2835 VSS nch l=0.04u w=0.8u
m5489 70912 4328 2831 VSS nch l=0.04u w=0.12u
m5490 70913 4328 2832 VSS nch l=0.04u w=0.12u
m5491 70914 2782 2836 VSS nch l=0.04u w=0.8u
m5492 70915 2786 2837 VSS nch l=0.04u w=0.8u
m5493 70916 2787 2838 VSS nch l=0.04u w=0.8u
m5494 70917 2788 2839 VSS nch l=0.04u w=0.8u
m5495 70918 2789 2840 VSS nch l=0.04u w=0.8u
m5496 70919 2790 2841 VSS nch l=0.04u w=0.8u
m5497 70920 2791 2842 VSS nch l=0.04u w=0.8u
m5498 70921 2792 2843 VSS nch l=0.04u w=0.8u
m5499 2850 155 VSS VSS nch l=0.04u w=0.4u
m5500 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5501 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5502 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5503 2844 2677 70902 VSS nch l=0.04u w=0.8u
m5504 2851 2813 VSS VSS nch l=0.04u w=0.4u
m5505 2852 2814 VSS VSS nch l=0.04u w=0.4u
m5506 VSS 2854 70903 VSS nch l=0.04u w=0.12u
m5507 VSS 2855 70904 VSS nch l=0.04u w=0.12u
m5508 VSS 2856 70905 VSS nch l=0.04u w=0.12u
m5509 VSS 2857 70906 VSS nch l=0.04u w=0.12u
m5510 VSS 2699 VSS VSS nch l=0.26u w=0.8u
m5511 VSS 2861 70908 VSS nch l=0.04u w=0.12u
m5512 VSS 2862 70909 VSS nch l=0.04u w=0.12u
m5513 70927 3228 2845 VSS nch l=0.04u w=0.8u
m5514 VSS 2678 70910 VSS nch l=0.04u w=0.8u
m5515 70928 3229 2846 VSS nch l=0.04u w=0.8u
m5516 VSS 2679 70911 VSS nch l=0.04u w=0.8u
m5517 VSS 2863 70912 VSS nch l=0.04u w=0.12u
m5518 VSS 2864 70913 VSS nch l=0.04u w=0.12u
m5519 70929 3230 2847 VSS nch l=0.04u w=0.8u
m5520 VSS 2680 70914 VSS nch l=0.04u w=0.8u
m5521 2853 4328 2833 VSS nch l=0.04u w=0.4u
m5522 VSS 2683 70915 VSS nch l=0.04u w=0.8u
m5523 VSS 2684 70916 VSS nch l=0.04u w=0.8u
m5524 70930 3231 2848 VSS nch l=0.04u w=0.8u
m5525 VSS 2685 70917 VSS nch l=0.04u w=0.8u
m5526 VSS 2686 70918 VSS nch l=0.04u w=0.8u
m5527 VSS 2687 70919 VSS nch l=0.04u w=0.8u
m5528 70931 3232 2849 VSS nch l=0.04u w=0.8u
m5529 VSS 2688 70920 VSS nch l=0.04u w=0.8u
m5530 VSS 2689 70921 VSS nch l=0.04u w=0.8u
m5531 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5532 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5533 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5534 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5535 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5536 2854 2825 VSS VSS nch l=0.04u w=0.4u
m5537 2855 2826 VSS VSS nch l=0.04u w=0.4u
m5538 2856 2827 VSS VSS nch l=0.04u w=0.4u
m5539 2857 2828 VSS VSS nch l=0.04u w=0.4u
m5540 2858 2859 VSS VSS nch l=0.04u w=0.8u
m5541 70938 2815 VSS VSS nch l=0.04u w=0.8u
m5542 2861 2829 VSS VSS nch l=0.04u w=0.4u
m5543 2862 2830 VSS VSS nch l=0.04u w=0.4u
m5544 70939 3500 70927 VSS nch l=0.04u w=0.8u
m5545 70940 3501 70928 VSS nch l=0.04u w=0.8u
m5546 2863 2831 VSS VSS nch l=0.04u w=0.4u
m5547 2864 2832 VSS VSS nch l=0.04u w=0.4u
m5548 70941 3502 70929 VSS nch l=0.04u w=0.8u
m5549 70942 2756 2853 VSS nch l=0.04u w=0.12u
m5550 70943 3503 70930 VSS nch l=0.04u w=0.8u
m5551 70944 3504 70931 VSS nch l=0.04u w=0.8u
m5552 70947 155 VSS VSS nch l=0.04u w=0.8u
m5553 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5554 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5555 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5556 2866 2739 VSS VSS nch l=0.04u w=0.4u
m5557 2860 2701 70938 VSS nch l=0.04u w=0.8u
m5558 VSS 3777 70939 VSS nch l=0.04u w=0.8u
m5559 VSS 3778 70940 VSS nch l=0.04u w=0.8u
m5560 VSS 3779 70941 VSS nch l=0.04u w=0.8u
m5561 2867 4328 VSS VSS nch l=0.04u w=0.4u
m5562 2868 4328 VSS VSS nch l=0.04u w=0.4u
m5563 VSS 2884 70942 VSS nch l=0.04u w=0.12u
m5564 VSS 3780 70943 VSS nch l=0.04u w=0.8u
m5565 VSS 3781 70944 VSS nch l=0.04u w=0.8u
m5566 70951 2834 VSS VSS nch l=0.04u w=0.8u
m5567 70952 2835 VSS VSS nch l=0.04u w=0.8u
m5568 70953 2836 VSS VSS nch l=0.04u w=0.8u
m5569 70954 2837 VSS VSS nch l=0.04u w=0.8u
m5570 70955 2838 VSS VSS nch l=0.04u w=0.8u
m5571 70956 2839 VSS VSS nch l=0.04u w=0.8u
m5572 70957 2840 VSS VSS nch l=0.04u w=0.8u
m5573 70958 2841 VSS VSS nch l=0.04u w=0.8u
m5574 70959 2842 VSS VSS nch l=0.04u w=0.8u
m5575 70960 2843 VSS VSS nch l=0.04u w=0.8u
m5576 2865 FBDIV[8] 70947 VSS nch l=0.04u w=0.8u
m5577 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5578 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5579 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5580 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5581 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5582 2879 2583 2866 VSS nch l=0.04u w=0.4u
m5583 2884 2853 VSS VSS nch l=0.04u w=0.4u
m5584 2885 4328 VSS VSS nch l=0.04u w=0.4u
m5585 2886 4328 VSS VSS nch l=0.04u w=0.4u
m5586 2887 4328 VSS VSS nch l=0.04u w=0.4u
m5587 2888 4328 VSS VSS nch l=0.04u w=0.4u
m5588 2880 4328 2861 VSS nch l=0.04u w=0.4u
m5589 2881 4328 2862 VSS nch l=0.04u w=0.4u
m5590 2869 2718 70951 VSS nch l=0.04u w=0.8u
m5591 2870 2723 70952 VSS nch l=0.04u w=0.8u
m5592 2882 4328 2863 VSS nch l=0.04u w=0.4u
m5593 2883 4328 2864 VSS nch l=0.04u w=0.4u
m5594 2871 2726 70953 VSS nch l=0.04u w=0.8u
m5595 2872 2727 70954 VSS nch l=0.04u w=0.8u
m5596 2873 2730 70955 VSS nch l=0.04u w=0.8u
m5597 2874 2731 70956 VSS nch l=0.04u w=0.8u
m5598 2875 2732 70957 VSS nch l=0.04u w=0.8u
m5599 2876 2735 70958 VSS nch l=0.04u w=0.8u
m5600 2877 2736 70959 VSS nch l=0.04u w=0.8u
m5601 2878 2737 70960 VSS nch l=0.04u w=0.8u
m5602 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5603 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5604 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5605 2583 2866 2879 VSS nch l=0.04u w=0.4u
m5606 2896 2926 VSS VSS nch l=0.04u w=0.4u
m5607 2897 2761 VSS VSS nch l=0.04u w=0.4u
m5608 70969 2809 2880 VSS nch l=0.04u w=0.12u
m5609 70970 2810 2881 VSS nch l=0.04u w=0.12u
m5610 VSS 2995 2889 VSS nch l=0.04u w=0.4u
m5611 VSS 2997 2890 VSS nch l=0.04u w=0.4u
m5612 70971 2811 2882 VSS nch l=0.04u w=0.12u
m5613 70972 2812 2883 VSS nch l=0.04u w=0.12u
m5614 VSS 3001 2891 VSS nch l=0.04u w=0.4u
m5615 2894 2867 2851 VSS nch l=0.04u w=0.4u
m5616 2895 2868 2852 VSS nch l=0.04u w=0.4u
m5617 VSS 3005 2892 VSS nch l=0.04u w=0.4u
m5618 VSS 3009 2893 VSS nch l=0.04u w=0.4u
m5619 VSS 2691 VSS VSS nch l=0.26u w=0.8u
m5620 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5621 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5622 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5623 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5624 70976 2850 VSS VSS nch l=0.04u w=0.8u
m5625 VSS 2926 2896 VSS nch l=0.04u w=0.4u
m5626 2906 2667 2897 VSS nch l=0.04u w=0.4u
m5627 VSS 2924 70969 VSS nch l=0.04u w=0.12u
m5628 VSS 2793 70970 VSS nch l=0.04u w=0.12u
m5629 VSS 2925 70971 VSS nch l=0.04u w=0.12u
m5630 VSS 2795 70972 VSS nch l=0.04u w=0.12u
m5631 70979 4328 2894 VSS nch l=0.04u w=0.12u
m5632 70980 4328 2895 VSS nch l=0.04u w=0.12u
m5633 2902 2885 2898 VSS nch l=0.04u w=0.4u
m5634 2903 2886 2899 VSS nch l=0.04u w=0.4u
m5635 2904 2887 2900 VSS nch l=0.04u w=0.4u
m5636 2905 2888 2798 VSS nch l=0.04u w=0.4u
m5637 2907 2908 VSS VSS nch l=0.04u w=0.8u
m5638 2910 2780 VSS VSS nch l=0.04u w=0.4u
m5639 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5640 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5641 2912 2781 VSS VSS nch l=0.04u w=0.4u
m5642 2914 2782 VSS VSS nch l=0.04u w=0.4u
m5643 2915 2786 VSS VSS nch l=0.04u w=0.4u
m5644 2916 2787 VSS VSS nch l=0.04u w=0.4u
m5645 2918 2788 VSS VSS nch l=0.04u w=0.4u
m5646 2919 2789 VSS VSS nch l=0.04u w=0.4u
m5647 2920 2790 VSS VSS nch l=0.04u w=0.4u
m5648 2922 2791 VSS VSS nch l=0.04u w=0.4u
m5649 2923 2792 VSS VSS nch l=0.04u w=0.4u
m5650 2901 2884 70976 VSS nch l=0.04u w=0.8u
m5651 VSS 2694 VSS VSS nch l=0.26u w=0.8u
m5652 2667 2897 2906 VSS nch l=0.04u w=0.4u
m5653 2924 2880 VSS VSS nch l=0.04u w=0.4u
m5654 2793 2881 VSS VSS nch l=0.04u w=0.4u
m5655 VSS 2706 VSS VSS nch l=0.26u w=0.8u
m5656 VSS 2707 VSS VSS nch l=0.26u w=0.8u
m5657 2925 2882 VSS VSS nch l=0.04u w=0.4u
m5658 2795 2883 VSS VSS nch l=0.04u w=0.4u
m5659 VSS 2710 VSS VSS nch l=0.26u w=0.8u
m5660 VSS 2711 VSS VSS nch l=0.26u w=0.8u
m5661 VSS 2944 70979 VSS nch l=0.04u w=0.12u
m5662 VSS 2945 70980 VSS nch l=0.04u w=0.12u
m5663 70993 4328 2902 VSS nch l=0.04u w=0.12u
m5664 70994 4328 2903 VSS nch l=0.04u w=0.12u
m5665 70995 4328 2904 VSS nch l=0.04u w=0.12u
m5666 70996 4328 2905 VSS nch l=0.04u w=0.12u
m5667 2927 2445 VSS VSS nch l=0.04u w=0.4u
m5668 2824 2678 2910 VSS nch l=0.04u w=0.4u
m5669 2929 2679 2912 VSS nch l=0.04u w=0.4u
m5670 2794 2680 2914 VSS nch l=0.04u w=0.4u
m5671 2774 2683 2915 VSS nch l=0.04u w=0.4u
m5672 2899 2684 2916 VSS nch l=0.04u w=0.4u
m5673 2931 2685 2918 VSS nch l=0.04u w=0.4u
m5674 2804 2686 2919 VSS nch l=0.04u w=0.4u
m5675 2798 2687 2920 VSS nch l=0.04u w=0.4u
m5676 2805 2688 2922 VSS nch l=0.04u w=0.4u
m5677 2808 2689 2923 VSS nch l=0.04u w=0.4u
m5678 2935 2934 VSS VSS nch l=0.04u w=0.8u
m5679 2936 2937 VSS VSS nch l=0.04u w=0.8u
m5680 2939 2938 VSS VSS nch l=0.04u w=0.8u
m5681 VSS 2720 VSS VSS nch l=0.26u w=0.8u
m5682 VSS 2721 VSS VSS nch l=0.26u w=0.8u
m5683 2940 2941 VSS VSS nch l=0.04u w=0.8u
m5684 2943 2942 VSS VSS nch l=0.04u w=0.8u
m5685 2944 2894 VSS VSS nch l=0.04u w=0.4u
m5686 2945 2895 VSS VSS nch l=0.04u w=0.4u
m5687 VSS 2960 70993 VSS nch l=0.04u w=0.12u
m5688 VSS 2961 70994 VSS nch l=0.04u w=0.12u
m5689 VSS 2962 70995 VSS nch l=0.04u w=0.12u
m5690 VSS 2963 70996 VSS nch l=0.04u w=0.12u
m5691 VSS 2977 2926 VSS nch l=0.04u w=0.4u
m5692 VSS 2879 2927 VSS nch l=0.04u w=0.4u
m5693 70999 2508 VSS VSS nch l=0.04u w=0.8u
m5694 2678 2910 2824 VSS nch l=0.04u w=0.4u
m5695 2679 2912 2929 VSS nch l=0.04u w=0.4u
m5696 2680 2914 2794 VSS nch l=0.04u w=0.4u
m5697 2683 2915 2774 VSS nch l=0.04u w=0.4u
m5698 2684 2916 2899 VSS nch l=0.04u w=0.4u
m5699 2685 2918 2931 VSS nch l=0.04u w=0.4u
m5700 2686 2919 2804 VSS nch l=0.04u w=0.4u
m5701 2687 2920 2798 VSS nch l=0.04u w=0.4u
m5702 2688 2922 2805 VSS nch l=0.04u w=0.4u
m5703 2689 2923 2808 VSS nch l=0.04u w=0.4u
m5704 VSS 2932 2932 VSS nch l=0.04u w=0.8u
m5705 2823 2964 2909 VSS nch l=0.04u w=0.4u
m5706 2928 2965 2911 VSS nch l=0.04u w=0.4u
m5707 2930 2966 2913 VSS nch l=0.04u w=0.4u
m5708 2743 2967 2917 VSS nch l=0.04u w=0.4u
m5709 2745 2968 2921 VSS nch l=0.04u w=0.4u
m5710 71000 2901 VSS VSS nch l=0.04u w=0.8u
m5711 71007 2896 VSS VSS nch l=0.04u w=0.8u
m5712 2956 2957 VSS VSS nch l=0.04u w=0.8u
m5713 2959 2958 VSS VSS nch l=0.04u w=0.8u
m5714 2960 2902 VSS VSS nch l=0.04u w=0.4u
m5715 2961 2903 VSS VSS nch l=0.04u w=0.4u
m5716 2962 2904 VSS VSS nch l=0.04u w=0.4u
m5717 2963 2905 VSS VSS nch l=0.04u w=0.4u
m5718 71008 2926 VSS VSS nch l=0.04u w=0.12u
m5719 2946 2465 70999 VSS nch l=0.04u w=0.8u
m5720 2964 2909 2823 VSS nch l=0.04u w=0.4u
m5721 2965 2911 2928 VSS nch l=0.04u w=0.4u
m5722 2966 2913 2930 VSS nch l=0.04u w=0.4u
m5723 2967 2917 2743 VSS nch l=0.04u w=0.4u
m5724 2968 2921 2745 VSS nch l=0.04u w=0.4u
m5725 2952 2865 71000 VSS nch l=0.04u w=0.8u
m5726 VSS 2954 2954 VSS nch l=0.04u w=0.8u
m5727 71025 3565 71007 VSS nch l=0.04u w=0.8u
m5728 2969 3013 VSS VSS nch l=0.04u w=0.4u
m5729 71026 2969 VSS VSS nch l=0.04u w=0.8u
m5730 2977 3085 71008 VSS nch l=0.04u w=0.12u
m5731 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m5732 2971 4328 2944 VSS nch l=0.04u w=0.4u
m5733 2972 4328 2945 VSS nch l=0.04u w=0.4u
m5734 71029 2445 VSS VSS nch l=0.04u w=0.8u
m5735 71030 110 VSS VSS nch l=0.04u w=0.8u
m5736 VSS 2947 2964 VSS nch l=0.04u w=0.4u
m5737 VSS 2948 2965 VSS nch l=0.04u w=0.4u
m5738 VSS 2949 2966 VSS nch l=0.04u w=0.4u
m5739 VSS 2950 2967 VSS nch l=0.04u w=0.4u
m5740 VSS 2951 2968 VSS nch l=0.04u w=0.4u
m5741 2955 4064 71025 VSS nch l=0.04u w=0.8u
m5742 VSS 3013 2969 VSS nch l=0.04u w=0.4u
m5743 71031 3484 71026 VSS nch l=0.04u w=0.8u
m5744 2993 4251 2977 VSS nch l=0.04u w=0.4u
m5745 VSS 2973 2973 VSS nch l=0.04u w=0.8u
m5746 VSS 2976 2976 VSS nch l=0.04u w=0.8u
m5747 71034 2867 2971 VSS nch l=0.04u w=0.12u
m5748 71035 2868 2972 VSS nch l=0.04u w=0.12u
m5749 2989 4328 2960 VSS nch l=0.04u w=0.4u
m5750 2990 4328 2961 VSS nch l=0.04u w=0.4u
m5751 2991 4328 2962 VSS nch l=0.04u w=0.4u
m5752 2992 4328 2963 VSS nch l=0.04u w=0.4u
m5753 2978 2465 71029 VSS nch l=0.04u w=0.8u
m5754 2994 2465 VSS VSS nch l=0.04u w=0.4u
m5755 2979 437 71030 VSS nch l=0.04u w=0.8u
m5756 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m5757 VSS 2980 2980 VSS nch l=0.04u w=0.8u
m5758 VSS 2983 2983 VSS nch l=0.04u w=0.8u
m5759 71036 3065 VSS VSS nch l=0.04u w=0.8u
m5760 71037 1877 VSS VSS nch l=0.04u w=0.8u
m5761 71038 2616 VSS VSS nch l=0.04u w=0.8u
m5762 71039 2616 VSS VSS nch l=0.04u w=0.8u
m5763 VSS 2984 2984 VSS nch l=0.04u w=0.8u
m5764 VSS 2987 2987 VSS nch l=0.04u w=0.8u
m5765 71040 FRAC[9] VSS VSS nch l=0.04u w=0.8u
m5766 VSS 3038 2988 VSS nch l=0.04u w=0.4u
m5767 71041 3066 VSS VSS nch l=0.04u w=0.8u
m5768 71042 3078 VSS VSS nch l=0.04u w=0.8u
m5769 71043 2900 VSS VSS nch l=0.04u w=0.8u
m5770 71044 2988 VSS VSS nch l=0.04u w=0.8u
m5771 71045 3079 VSS VSS nch l=0.04u w=0.8u
m5772 71046 FRAC[9] VSS VSS nch l=0.04u w=0.8u
m5773 71047 2988 VSS VSS nch l=0.04u w=0.8u
m5774 3012 3062 VSS VSS nch l=0.04u w=0.4u
m5775 2970 3953 71031 VSS nch l=0.04u w=0.8u
m5776 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m5777 VSS 1146 71034 VSS nch l=0.04u w=0.12u
m5778 VSS 3018 71035 VSS nch l=0.04u w=0.12u
m5779 71049 2885 2989 VSS nch l=0.04u w=0.12u
m5780 71050 2886 2990 VSS nch l=0.04u w=0.12u
m5781 71051 2887 2991 VSS nch l=0.04u w=0.12u
m5782 71052 2888 2992 VSS nch l=0.04u w=0.12u
m5783 3016 2508 2994 VSS nch l=0.04u w=0.4u
m5784 71053 3144 2995 VSS nch l=0.04u w=0.8u
m5785 2996 3063 71036 VSS nch l=0.04u w=0.8u
m5786 71054 3146 2997 VSS nch l=0.04u w=0.8u
m5787 2998 3064 71037 VSS nch l=0.04u w=0.8u
m5788 2999 3206 71038 VSS nch l=0.04u w=0.8u
m5789 3000 3207 71039 VSS nch l=0.04u w=0.8u
m5790 71055 3148 3001 VSS nch l=0.04u w=0.8u
m5791 3002 3065 71040 VSS nch l=0.04u w=0.8u
m5792 3003 131 71041 VSS nch l=0.04u w=0.8u
m5793 3004 3066 71042 VSS nch l=0.04u w=0.8u
m5794 71056 3152 3005 VSS nch l=0.04u w=0.8u
m5795 3006 3023 71043 VSS nch l=0.04u w=0.8u
m5796 3007 3067 71044 VSS nch l=0.04u w=0.8u
m5797 3008 3068 71045 VSS nch l=0.04u w=0.8u
m5798 71057 3156 3009 VSS nch l=0.04u w=0.8u
m5799 3010 3024 71046 VSS nch l=0.04u w=0.8u
m5800 3011 FBDIV[9] 71047 VSS nch l=0.04u w=0.8u
m5801 VSS 3062 3012 VSS nch l=0.04u w=0.4u
m5802 3017 2955 VSS VSS nch l=0.04u w=0.4u
m5803 VSS 3041 3013 VSS nch l=0.04u w=0.4u
m5804 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m5805 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m5806 VSS 3015 3015 VSS nch l=0.04u w=0.8u
m5807 1146 2971 VSS VSS nch l=0.04u w=0.4u
m5808 3018 2972 VSS VSS nch l=0.04u w=0.4u
m5809 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m5810 VSS 3023 71049 VSS nch l=0.04u w=0.12u
m5811 VSS 2796 71050 VSS nch l=0.04u w=0.12u
m5812 VSS 3024 71051 VSS nch l=0.04u w=0.12u
m5813 VSS 2799 71052 VSS nch l=0.04u w=0.12u
m5814 VSS 3044 2993 VSS nch l=0.04u w=0.4u
m5815 2508 2994 3016 VSS nch l=0.04u w=0.4u
m5816 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m5817 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m5818 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m5819 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m5820 3019 2978 VSS VSS nch l=0.04u w=0.4u
m5821 3020 437 VSS VSS nch l=0.04u w=0.4u
m5822 VSS 3046 71053 VSS nch l=0.04u w=0.8u
m5823 VSS 3048 71054 VSS nch l=0.04u w=0.8u
m5824 VSS 3050 71055 VSS nch l=0.04u w=0.8u
m5825 VSS 3055 71056 VSS nch l=0.04u w=0.8u
m5826 VSS 3059 71057 VSS nch l=0.04u w=0.8u
m5827 3012 3062 VSS VSS nch l=0.04u w=0.4u
m5828 3021 4328 VSS VSS nch l=0.04u w=0.4u
m5829 71060 3013 VSS VSS nch l=0.04u w=0.12u
m5830 3022 2970 VSS VSS nch l=0.04u w=0.4u
m5831 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m5832 3023 2989 VSS VSS nch l=0.04u w=0.4u
m5833 2796 2990 VSS VSS nch l=0.04u w=0.4u
m5834 3024 2991 VSS VSS nch l=0.04u w=0.4u
m5835 2799 2992 VSS VSS nch l=0.04u w=0.4u
m5836 71061 2993 VSS VSS nch l=0.04u w=0.12u
m5837 3025 110 3020 VSS nch l=0.04u w=0.4u
m5838 VSS 3062 3012 VSS nch l=0.04u w=0.4u
m5839 3026 3063 VSS VSS nch l=0.04u w=0.4u
m5840 3027 3064 VSS VSS nch l=0.04u w=0.4u
m5841 3028 2999 VSS VSS nch l=0.04u w=0.4u
m5842 3029 3000 VSS VSS nch l=0.04u w=0.4u
m5843 3030 3065 VSS VSS nch l=0.04u w=0.4u
m5844 3031 131 VSS VSS nch l=0.04u w=0.4u
m5845 3032 3066 VSS VSS nch l=0.04u w=0.4u
m5846 3033 3023 VSS VSS nch l=0.04u w=0.4u
m5847 3034 3067 VSS VSS nch l=0.04u w=0.4u
m5848 3035 3068 VSS VSS nch l=0.04u w=0.4u
m5849 3036 3024 VSS VSS nch l=0.04u w=0.4u
m5850 3037 FBDIV[9] VSS VSS nch l=0.04u w=0.4u
m5851 71063 3017 VSS VSS nch l=0.04u w=0.8u
m5852 3041 3141 71060 VSS nch l=0.04u w=0.12u
m5853 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m5854 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m5855 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m5856 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m5857 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m5858 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m5859 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m5860 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m5861 3044 4251 71061 VSS nch l=0.04u w=0.12u
m5862 3042 912 VSS VSS nch l=0.04u w=0.4u
m5863 3043 4328 VSS VSS nch l=0.04u w=0.4u
m5864 110 3020 3025 VSS nch l=0.04u w=0.4u
m5865 71064 2909 VSS VSS nch l=0.04u w=0.8u
m5866 3047 3065 3026 VSS nch l=0.04u w=0.4u
m5867 71065 2911 VSS VSS nch l=0.04u w=0.8u
m5868 3049 1877 3027 VSS nch l=0.04u w=0.4u
m5869 71066 2913 VSS VSS nch l=0.04u w=0.8u
m5870 3051 FRAC[9] 3030 VSS nch l=0.04u w=0.4u
m5871 3053 3066 3031 VSS nch l=0.04u w=0.4u
m5872 3054 3078 3032 VSS nch l=0.04u w=0.4u
m5873 71067 2917 VSS VSS nch l=0.04u w=0.8u
m5874 3056 2900 3033 VSS nch l=0.04u w=0.4u
m5875 3057 2988 3034 VSS nch l=0.04u w=0.4u
m5876 3058 3079 3035 VSS nch l=0.04u w=0.4u
m5877 71068 2921 VSS VSS nch l=0.04u w=0.8u
m5878 3060 FRAC[9] 3036 VSS nch l=0.04u w=0.4u
m5879 3061 2988 3037 VSS nch l=0.04u w=0.4u
m5880 3052 3021 3038 VSS nch l=0.04u w=0.4u
m5881 71069 4351 71063 VSS nch l=0.04u w=0.8u
m5882 3069 4251 3041 VSS nch l=0.04u w=0.4u
m5883 3040 3070 2970 VSS nch l=0.04u w=0.4u
m5884 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m5885 3071 3085 3044 VSS nch l=0.04u w=0.4u
m5886 3072 1146 3042 VSS nch l=0.04u w=0.4u
m5887 3073 4328 VSS VSS nch l=0.04u w=0.4u
m5888 3074 4328 VSS VSS nch l=0.04u w=0.4u
m5889 3075 4328 VSS VSS nch l=0.04u w=0.4u
m5890 3076 4328 VSS VSS nch l=0.04u w=0.4u
m5891 71070 3016 3045 VSS nch l=0.04u w=0.8u
m5892 3046 2947 71064 VSS nch l=0.04u w=0.8u
m5893 3065 3026 3047 VSS nch l=0.04u w=0.4u
m5894 3048 2948 71065 VSS nch l=0.04u w=0.8u
m5895 1877 3027 3049 VSS nch l=0.04u w=0.4u
m5896 3050 2949 71066 VSS nch l=0.04u w=0.8u
m5897 FRAC[9] 3030 3051 VSS nch l=0.04u w=0.4u
m5898 3066 3031 3053 VSS nch l=0.04u w=0.4u
m5899 3078 3032 3054 VSS nch l=0.04u w=0.4u
m5900 3055 2950 71067 VSS nch l=0.04u w=0.8u
m5901 2900 3033 3056 VSS nch l=0.04u w=0.4u
m5902 2988 3034 3057 VSS nch l=0.04u w=0.4u
m5903 3079 3035 3058 VSS nch l=0.04u w=0.4u
m5904 3059 2951 71068 VSS nch l=0.04u w=0.8u
m5905 FRAC[9] 3036 3060 VSS nch l=0.04u w=0.4u
m5906 2988 3037 3061 VSS nch l=0.04u w=0.4u
m5907 VSS 4062 3062 VSS nch l=0.04u w=0.4u
m5908 3080 4328 VSS VSS nch l=0.04u w=0.4u
m5909 3081 4328 VSS VSS nch l=0.04u w=0.4u
m5910 3082 4328 VSS VSS nch l=0.04u w=0.4u
m5911 3083 4328 VSS VSS nch l=0.04u w=0.4u
m5912 71071 4328 3052 VSS nch l=0.04u w=0.12u
m5913 3039 3484 71069 VSS nch l=0.04u w=0.8u
m5914 3070 2970 3040 VSS nch l=0.04u w=0.4u
m5915 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m5916 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m5917 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m5918 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m5919 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m5920 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m5921 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m5922 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m5923 1146 3042 3072 VSS nch l=0.04u w=0.4u
m5924 3084 3043 3018 VSS nch l=0.04u w=0.4u
m5925 VSS 2844 71070 VSS nch l=0.04u w=0.8u
m5926 VSS 3101 71071 VSS nch l=0.04u w=0.12u
m5927 VSS 3118 3069 VSS nch l=0.04u w=0.4u
m5928 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m5929 VSS 4251 3085 VSS nch l=0.04u w=0.4u
m5930 71088 4328 3084 VSS nch l=0.04u w=0.12u
m5931 3092 3073 3086 VSS nch l=0.04u w=0.4u
m5932 3093 3074 2931 VSS nch l=0.04u w=0.4u
m5933 3094 3075 3087 VSS nch l=0.04u w=0.4u
m5934 3095 3076 2805 VSS nch l=0.04u w=0.4u
m5935 2630 3096 VSS VSS nch l=0.04u w=0.8u
m5936 71089 3025 3088 VSS nch l=0.04u w=0.8u
m5937 3101 3052 VSS VSS nch l=0.04u w=0.4u
m5938 3102 3117 VSS VSS nch l=0.04u w=0.4u
m5939 3097 3080 3090 VSS nch l=0.04u w=0.4u
m5940 3098 3081 3091 VSS nch l=0.04u w=0.4u
m5941 3099 3082 3028 VSS nch l=0.04u w=0.4u
m5942 3100 3083 3029 VSS nch l=0.04u w=0.4u
m5943 3113 3039 VSS VSS nch l=0.04u w=0.4u
m5944 71090 3069 VSS VSS nch l=0.04u w=0.12u
m5945 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m5946 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m5947 3114 4062 VSS VSS nch l=0.04u w=0.4u
m5948 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m5949 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m5950 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m5951 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m5952 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m5953 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m5954 VSS 3119 71088 VSS nch l=0.04u w=0.12u
m5955 71091 4328 3092 VSS nch l=0.04u w=0.12u
m5956 71092 4328 3093 VSS nch l=0.04u w=0.12u
m5957 71093 4328 3094 VSS nch l=0.04u w=0.12u
m5958 71094 4328 3095 VSS nch l=0.04u w=0.12u
m5959 71095 3045 VSS VSS nch l=0.04u w=0.8u
m5960 VSS 2860 71089 VSS nch l=0.04u w=0.8u
m5961 71096 4328 3097 VSS nch l=0.04u w=0.12u
m5962 71097 4328 3098 VSS nch l=0.04u w=0.12u
m5963 2947 3123 2925 VSS nch l=0.04u w=0.4u
m5964 71098 3047 3103 VSS nch l=0.04u w=0.8u
m5965 2948 3124 2054 VSS nch l=0.04u w=0.4u
m5966 71099 3049 3104 VSS nch l=0.04u w=0.8u
m5967 71100 4328 3099 VSS nch l=0.04u w=0.12u
m5968 71101 4328 3100 VSS nch l=0.04u w=0.12u
m5969 2949 3125 FRAC[15] VSS nch l=0.04u w=0.4u
m5970 71102 3051 3105 VSS nch l=0.04u w=0.8u
m5971 71103 3053 3106 VSS nch l=0.04u w=0.8u
m5972 71104 3054 3107 VSS nch l=0.04u w=0.8u
m5973 2950 3126 2745 VSS nch l=0.04u w=0.4u
m5974 71105 3056 3108 VSS nch l=0.04u w=0.8u
m5975 71106 3057 3109 VSS nch l=0.04u w=0.8u
m5976 71107 3058 3110 VSS nch l=0.04u w=0.8u
m5977 2951 3127 FRAC[15] VSS nch l=0.04u w=0.4u
m5978 71108 3060 3111 VSS nch l=0.04u w=0.8u
m5979 71109 3061 3112 VSS nch l=0.04u w=0.8u
m5980 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m5981 3118 4251 71090 VSS nch l=0.04u w=0.12u
m5982 3119 3084 VSS VSS nch l=0.04u w=0.4u
m5983 VSS 3132 71091 VSS nch l=0.04u w=0.12u
m5984 VSS 3133 71092 VSS nch l=0.04u w=0.12u
m5985 VSS 3134 71093 VSS nch l=0.04u w=0.12u
m5986 VSS 3135 71094 VSS nch l=0.04u w=0.12u
m5987 71110 3173 VSS VSS nch l=0.04u w=0.8u
m5988 3120 3120 VSS VSS nch l=0.04u w=0.8u
m5989 3115 2946 71095 VSS nch l=0.04u w=0.8u
m5990 VSS 3137 71096 VSS nch l=0.04u w=0.12u
m5991 VSS 3138 71097 VSS nch l=0.04u w=0.12u
m5992 3123 2925 2947 VSS nch l=0.04u w=0.4u
m5993 VSS 2869 71098 VSS nch l=0.04u w=0.8u
m5994 3124 2054 2948 VSS nch l=0.04u w=0.4u
m5995 VSS 2870 71099 VSS nch l=0.04u w=0.8u
m5996 VSS 3139 71100 VSS nch l=0.04u w=0.12u
m5997 VSS 3140 71101 VSS nch l=0.04u w=0.12u
m5998 3125 FRAC[15] 2949 VSS nch l=0.04u w=0.4u
m5999 VSS 2871 71102 VSS nch l=0.04u w=0.8u
m6000 3121 4328 3101 VSS nch l=0.04u w=0.4u
m6001 VSS 2872 71103 VSS nch l=0.04u w=0.8u
m6002 VSS 2873 71104 VSS nch l=0.04u w=0.8u
m6003 3126 2745 2950 VSS nch l=0.04u w=0.4u
m6004 VSS 2874 71105 VSS nch l=0.04u w=0.8u
m6005 VSS 2875 71106 VSS nch l=0.04u w=0.8u
m6006 VSS 2876 71107 VSS nch l=0.04u w=0.8u
m6007 3127 FRAC[15] 2951 VSS nch l=0.04u w=0.4u
m6008 VSS 2877 71108 VSS nch l=0.04u w=0.8u
m6009 VSS 2878 71109 VSS nch l=0.04u w=0.8u
m6010 3116 3122 3117 VSS nch l=0.04u w=0.4u
m6011 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m6012 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m6013 3128 3141 3118 VSS nch l=0.04u w=0.4u
m6014 71111 3113 VSS VSS nch l=0.04u w=0.8u
m6015 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m6016 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m6017 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m6018 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m6019 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m6020 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m6021 71112 4062 VSS VSS nch l=0.04u w=0.8u
m6022 3131 4328 VSS VSS nch l=0.04u w=0.4u
m6023 3132 3092 VSS VSS nch l=0.04u w=0.4u
m6024 3133 3093 VSS VSS nch l=0.04u w=0.4u
m6025 3134 3094 VSS VSS nch l=0.04u w=0.4u
m6026 3135 3095 VSS VSS nch l=0.04u w=0.4u
m6027 3071 3218 71110 VSS nch l=0.04u w=0.8u
m6028 71113 3088 VSS VSS nch l=0.04u w=0.8u
m6029 3137 3097 VSS VSS nch l=0.04u w=0.4u
m6030 3138 3098 VSS VSS nch l=0.04u w=0.4u
m6031 VSS 2924 3123 VSS nch l=0.04u w=0.4u
m6032 VSS 2930 3124 VSS nch l=0.04u w=0.4u
m6033 3139 3099 VSS VSS nch l=0.04u w=0.4u
m6034 3140 3100 VSS VSS nch l=0.04u w=0.4u
m6035 VSS 2925 3125 VSS nch l=0.04u w=0.4u
m6036 71114 3021 3121 VSS nch l=0.04u w=0.12u
m6037 VSS 2855 3126 VSS nch l=0.04u w=0.4u
m6038 VSS 2857 3127 VSS nch l=0.04u w=0.4u
m6039 3122 3117 3116 VSS nch l=0.04u w=0.4u
m6040 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m6041 3129 3953 71111 VSS nch l=0.04u w=0.8u
m6042 3130 1962 71112 VSS nch l=0.04u w=0.8u
m6043 71115 3218 3071 VSS nch l=0.04u w=0.8u
m6044 3142 4328 3119 VSS nch l=0.04u w=0.4u
m6045 3143 3016 VSS VSS nch l=0.04u w=0.4u
m6046 3136 2979 71113 VSS nch l=0.04u w=0.8u
m6047 VSS 3169 71114 VSS nch l=0.04u w=0.12u
m6048 71116 3103 VSS VSS nch l=0.04u w=0.8u
m6049 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m6050 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m6051 71117 3104 VSS VSS nch l=0.04u w=0.8u
m6052 71118 3105 VSS VSS nch l=0.04u w=0.8u
m6053 71119 3106 VSS VSS nch l=0.04u w=0.8u
m6054 71120 3107 VSS VSS nch l=0.04u w=0.8u
m6055 71121 3108 VSS VSS nch l=0.04u w=0.8u
m6056 71122 3109 VSS VSS nch l=0.04u w=0.8u
m6057 71123 3110 VSS VSS nch l=0.04u w=0.8u
m6058 71124 3111 VSS VSS nch l=0.04u w=0.8u
m6059 71125 3112 VSS VSS nch l=0.04u w=0.8u
m6060 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m6061 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m6062 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m6063 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m6064 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m6065 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m6066 VSS 4251 3141 VSS nch l=0.04u w=0.4u
m6067 3159 3131 3072 VSS nch l=0.04u w=0.4u
m6068 VSS 3173 71115 VSS nch l=0.04u w=0.8u
m6069 71126 3043 3142 VSS nch l=0.04u w=0.12u
m6070 3160 4328 3132 VSS nch l=0.04u w=0.4u
m6071 3161 4328 3133 VSS nch l=0.04u w=0.4u
m6072 3162 4328 3134 VSS nch l=0.04u w=0.4u
m6073 3163 4328 3135 VSS nch l=0.04u w=0.4u
m6074 VSS 2933 VSS VSS nch l=0.26u w=0.8u
m6075 3164 2844 3143 VSS nch l=0.04u w=0.4u
m6076 3169 3121 VSS VSS nch l=0.04u w=0.4u
m6077 3165 4328 3137 VSS nch l=0.04u w=0.4u
m6078 3166 4328 3138 VSS nch l=0.04u w=0.4u
m6079 71127 2924 3144 VSS nch l=0.04u w=0.8u
m6080 3145 2996 71116 VSS nch l=0.04u w=0.8u
m6081 71128 2930 3146 VSS nch l=0.04u w=0.8u
m6082 3147 2998 71117 VSS nch l=0.04u w=0.8u
m6083 3167 4328 3139 VSS nch l=0.04u w=0.4u
m6084 3168 4328 3140 VSS nch l=0.04u w=0.4u
m6085 71129 2925 3148 VSS nch l=0.04u w=0.8u
m6086 3149 3002 71118 VSS nch l=0.04u w=0.8u
m6087 3150 3003 71119 VSS nch l=0.04u w=0.8u
m6088 3151 3004 71120 VSS nch l=0.04u w=0.8u
m6089 71130 2855 3152 VSS nch l=0.04u w=0.8u
m6090 3153 3006 71121 VSS nch l=0.04u w=0.8u
m6091 3154 3007 71122 VSS nch l=0.04u w=0.8u
m6092 3155 3008 71123 VSS nch l=0.04u w=0.8u
m6093 71131 2857 3156 VSS nch l=0.04u w=0.8u
m6094 3157 3010 71124 VSS nch l=0.04u w=0.8u
m6095 3158 3011 71125 VSS nch l=0.04u w=0.8u
m6096 3170 4062 VSS VSS nch l=0.04u w=0.4u
m6097 3171 3129 VSS VSS nch l=0.04u w=0.4u
m6098 71132 3114 VSS VSS nch l=0.04u w=0.8u
m6099 71133 4328 3159 VSS nch l=0.04u w=0.12u
m6100 VSS 61 71126 VSS nch l=0.04u w=0.12u
m6101 71134 3073 3160 VSS nch l=0.04u w=0.12u
m6102 71135 3074 3161 VSS nch l=0.04u w=0.12u
m6103 71136 3075 3162 VSS nch l=0.04u w=0.12u
m6104 71137 3076 3163 VSS nch l=0.04u w=0.12u
m6105 3174 3175 VSS VSS nch l=0.04u w=0.8u
m6106 2844 3143 3164 VSS nch l=0.04u w=0.4u
m6107 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m6108 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m6109 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m6110 3176 3025 VSS VSS nch l=0.04u w=0.4u
m6111 71138 3080 3165 VSS nch l=0.04u w=0.12u
m6112 71139 3081 3166 VSS nch l=0.04u w=0.12u
m6113 VSS 2925 71127 VSS nch l=0.04u w=0.8u
m6114 VSS 2054 71128 VSS nch l=0.04u w=0.8u
m6115 71140 3082 3167 VSS nch l=0.04u w=0.12u
m6116 71141 3083 3168 VSS nch l=0.04u w=0.12u
m6117 VSS FRAC[15] 71129 VSS nch l=0.04u w=0.8u
m6118 VSS 2953 VSS VSS nch l=0.26u w=0.8u
m6119 VSS 2745 71130 VSS nch l=0.04u w=0.8u
m6120 VSS FRAC[15] 71131 VSS nch l=0.04u w=0.8u
m6121 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m6122 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m6123 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m6124 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m6125 71143 3249 VSS VSS nch l=0.04u w=0.8u
m6126 3172 3040 71132 VSS nch l=0.04u w=0.8u
m6127 VSS 3200 71133 VSS nch l=0.04u w=0.12u
m6128 61 3142 VSS VSS nch l=0.04u w=0.4u
m6129 VSS 3201 71134 VSS nch l=0.04u w=0.12u
m6130 VSS 2797 71135 VSS nch l=0.04u w=0.12u
m6131 VSS 3202 71136 VSS nch l=0.04u w=0.12u
m6132 VSS 2800 71137 VSS nch l=0.04u w=0.12u
m6133 71144 3301 3173 VSS nch l=0.04u w=0.8u
m6134 3180 2860 3176 VSS nch l=0.04u w=0.4u
m6135 VSS 3203 71138 VSS nch l=0.04u w=0.12u
m6136 VSS 3063 71139 VSS nch l=0.04u w=0.12u
m6137 VSS 3204 71140 VSS nch l=0.04u w=0.12u
m6138 VSS 3065 71141 VSS nch l=0.04u w=0.12u
m6139 3182 3181 VSS VSS nch l=0.04u w=0.8u
m6140 3184 3047 VSS VSS nch l=0.04u w=0.4u
m6141 3186 3049 VSS VSS nch l=0.04u w=0.4u
m6142 3188 3051 VSS VSS nch l=0.04u w=0.4u
m6143 3189 3053 VSS VSS nch l=0.04u w=0.4u
m6144 3190 3054 VSS VSS nch l=0.04u w=0.4u
m6145 3192 3056 VSS VSS nch l=0.04u w=0.4u
m6146 3193 3057 VSS VSS nch l=0.04u w=0.4u
m6147 3194 3058 VSS VSS nch l=0.04u w=0.4u
m6148 3196 3060 VSS VSS nch l=0.04u w=0.4u
m6149 3197 3061 VSS VSS nch l=0.04u w=0.4u
m6150 71146 4062 VSS VSS nch l=0.04u w=0.8u
m6151 3128 3290 71143 VSS nch l=0.04u w=0.8u
m6152 3177 3199 3129 VSS nch l=0.04u w=0.4u
m6153 3200 3159 VSS VSS nch l=0.04u w=0.4u
m6154 3201 3160 VSS VSS nch l=0.04u w=0.4u
m6155 2797 3161 VSS VSS nch l=0.04u w=0.4u
m6156 3202 3162 VSS VSS nch l=0.04u w=0.4u
m6157 2800 3163 VSS VSS nch l=0.04u w=0.4u
m6158 VSS 3272 71144 VSS nch l=0.04u w=0.8u
m6159 VSS 2974 VSS VSS nch l=0.26u w=0.8u
m6160 VSS 2975 VSS VSS nch l=0.26u w=0.8u
m6161 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m6162 VSS 3178 3178 VSS nch l=0.04u w=0.8u
m6163 2860 3176 3180 VSS nch l=0.04u w=0.4u
m6164 3203 3165 VSS VSS nch l=0.04u w=0.4u
m6165 3063 3166 VSS VSS nch l=0.04u w=0.4u
m6166 VSS 2981 VSS VSS nch l=0.26u w=0.8u
m6167 VSS 2982 VSS VSS nch l=0.26u w=0.8u
m6168 3204 3167 VSS VSS nch l=0.04u w=0.4u
m6169 3065 3168 VSS VSS nch l=0.04u w=0.4u
m6170 VSS 2985 VSS VSS nch l=0.26u w=0.8u
m6171 VSS 2986 VSS VSS nch l=0.26u w=0.8u
m6172 3205 2445 VSS VSS nch l=0.04u w=0.4u
m6173 3091 2869 3184 VSS nch l=0.04u w=0.4u
m6174 3207 2870 3186 VSS nch l=0.04u w=0.4u
m6175 3064 2871 3188 VSS nch l=0.04u w=0.4u
m6176 3038 2872 3189 VSS nch l=0.04u w=0.4u
m6177 3211 2873 3190 VSS nch l=0.04u w=0.4u
m6178 2898 2874 3192 VSS nch l=0.04u w=0.4u
m6179 3078 2875 3193 VSS nch l=0.04u w=0.4u
m6180 3067 2876 3194 VSS nch l=0.04u w=0.4u
m6181 2900 2877 3196 VSS nch l=0.04u w=0.4u
m6182 3079 2878 3197 VSS nch l=0.04u w=0.4u
m6183 3198 320 71146 VSS nch l=0.04u w=0.8u
m6184 71154 3290 3128 VSS nch l=0.04u w=0.8u
m6185 3199 3129 3177 VSS nch l=0.04u w=0.4u
m6186 71155 3172 VSS VSS nch l=0.04u w=0.8u
m6187 3213 3214 VSS VSS nch l=0.04u w=0.8u
m6188 3216 3215 VSS VSS nch l=0.04u w=0.8u
m6189 3217 2098 VSS VSS nch l=0.04u w=0.4u
m6190 3219 3220 VSS VSS nch l=0.04u w=0.8u
m6191 3222 3221 VSS VSS nch l=0.04u w=0.8u
m6192 3223 3224 VSS VSS nch l=0.04u w=0.8u
m6193 3226 3225 VSS VSS nch l=0.04u w=0.8u
m6194 VSS 3164 3205 VSS nch l=0.04u w=0.4u
m6195 71157 2508 VSS VSS nch l=0.04u w=0.8u
m6196 2869 3184 3091 VSS nch l=0.04u w=0.4u
m6197 2870 3186 3207 VSS nch l=0.04u w=0.4u
m6198 2871 3188 3064 VSS nch l=0.04u w=0.4u
m6199 VSS 3210 3210 VSS nch l=0.04u w=0.8u
m6200 2872 3189 3038 VSS nch l=0.04u w=0.4u
m6201 2873 3190 3211 VSS nch l=0.04u w=0.4u
m6202 2874 3192 2898 VSS nch l=0.04u w=0.4u
m6203 2875 3193 3078 VSS nch l=0.04u w=0.4u
m6204 2876 3194 3067 VSS nch l=0.04u w=0.4u
m6205 2877 3196 2900 VSS nch l=0.04u w=0.4u
m6206 2878 3197 3079 VSS nch l=0.04u w=0.4u
m6207 3090 3243 3183 VSS nch l=0.04u w=0.4u
m6208 3206 3244 3185 VSS nch l=0.04u w=0.4u
m6209 3208 3245 3187 VSS nch l=0.04u w=0.4u
m6210 2742 3246 3191 VSS nch l=0.04u w=0.4u
m6211 2744 3247 3195 VSS nch l=0.04u w=0.4u
m6212 VSS 3249 71154 VSS nch l=0.04u w=0.8u
m6213 3212 3130 71155 VSS nch l=0.04u w=0.8u
m6214 3233 4328 3200 VSS nch l=0.04u w=0.4u
m6215 VSS 3014 VSS VSS nch l=0.26u w=0.8u
m6216 3234 3018 3217 VSS nch l=0.04u w=0.4u
m6217 3235 4328 VSS VSS nch l=0.04u w=0.4u
m6218 3236 4328 VSS VSS nch l=0.04u w=0.4u
m6219 3237 4328 VSS VSS nch l=0.04u w=0.4u
m6220 3238 4328 VSS VSS nch l=0.04u w=0.4u
m6221 71163 FBDIV[10] 3218 VSS nch l=0.04u w=0.8u
m6222 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6223 3227 2906 71157 VSS nch l=0.04u w=0.8u
m6224 3243 3183 3090 VSS nch l=0.04u w=0.4u
m6225 3244 3185 3206 VSS nch l=0.04u w=0.4u
m6226 3245 3187 3208 VSS nch l=0.04u w=0.4u
m6227 3246 3191 2742 VSS nch l=0.04u w=0.4u
m6228 3247 3195 2744 VSS nch l=0.04u w=0.4u
m6229 71165 3170 VSS VSS nch l=0.04u w=0.8u
m6230 3250 4062 VSS VSS nch l=0.04u w=0.4u
m6231 71182 3130 3212 VSS nch l=0.04u w=0.8u
m6232 71184 3131 3233 VSS nch l=0.04u w=0.12u
m6233 3252 3251 VSS VSS nch l=0.04u w=0.8u
m6234 3018 3217 3234 VSS nch l=0.04u w=0.4u
m6235 VSS 4062 71163 VSS nch l=0.04u w=0.8u
m6236 VSS 3239 3239 VSS nch l=0.04u w=0.8u
m6237 VSS 3242 3242 VSS nch l=0.04u w=0.8u
m6238 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6239 71187 2445 VSS VSS nch l=0.04u w=0.8u
m6240 71188 110 VSS VSS nch l=0.04u w=0.8u
m6241 VSS 3228 3243 VSS nch l=0.04u w=0.4u
m6242 VSS 3229 3244 VSS nch l=0.04u w=0.4u
m6243 VSS 3230 3245 VSS nch l=0.04u w=0.4u
m6244 VSS 3231 3246 VSS nch l=0.04u w=0.4u
m6245 VSS 3232 3247 VSS nch l=0.04u w=0.4u
m6246 3248 3116 71165 VSS nch l=0.04u w=0.8u
m6247 71189 3381 3249 VSS nch l=0.04u w=0.8u
m6248 VSS 3172 71182 VSS nch l=0.04u w=0.8u
m6249 VSS 3287 71184 VSS nch l=0.04u w=0.12u
m6250 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6251 3266 3235 3253 VSS nch l=0.04u w=0.4u
m6252 3267 3236 3211 VSS nch l=0.04u w=0.4u
m6253 3268 3237 3254 VSS nch l=0.04u w=0.4u
m6254 3269 3238 3067 VSS nch l=0.04u w=0.4u
m6255 3255 2906 71187 VSS nch l=0.04u w=0.8u
m6256 3273 2906 VSS VSS nch l=0.04u w=0.4u
m6257 3256 731 71188 VSS nch l=0.04u w=0.8u
m6258 VSS 3257 3257 VSS nch l=0.04u w=0.8u
m6259 VSS 3260 3260 VSS nch l=0.04u w=0.8u
m6260 71193 3338 VSS VSS nch l=0.04u w=0.8u
m6261 71194 1908 VSS VSS nch l=0.04u w=0.8u
m6262 71195 2616 VSS VSS nch l=0.04u w=0.8u
m6263 71196 2616 VSS VSS nch l=0.04u w=0.8u
m6264 VSS 3261 3261 VSS nch l=0.04u w=0.8u
m6265 VSS 3264 3264 VSS nch l=0.04u w=0.8u
m6266 71197 FRAC[10] VSS VSS nch l=0.04u w=0.8u
m6267 VSS 3315 3265 VSS nch l=0.04u w=0.4u
m6268 71198 3339 VSS VSS nch l=0.04u w=0.8u
m6269 71199 3352 VSS VSS nch l=0.04u w=0.8u
m6270 71200 3254 VSS VSS nch l=0.04u w=0.8u
m6271 71201 3265 VSS VSS nch l=0.04u w=0.8u
m6272 71202 3353 VSS VSS nch l=0.04u w=0.8u
m6273 71203 FRAC[10] VSS VSS nch l=0.04u w=0.8u
m6274 71204 3265 VSS VSS nch l=0.04u w=0.8u
m6275 VSS 3344 71189 VSS nch l=0.04u w=0.8u
m6276 71205 4062 VSS VSS nch l=0.04u w=0.8u
m6277 3287 3233 VSS VSS nch l=0.04u w=0.4u
m6278 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6279 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6280 VSS 3271 3271 VSS nch l=0.04u w=0.8u
m6281 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6282 71206 4328 3266 VSS nch l=0.04u w=0.12u
m6283 71207 4328 3267 VSS nch l=0.04u w=0.12u
m6284 71208 4328 3268 VSS nch l=0.04u w=0.12u
m6285 71209 4328 3269 VSS nch l=0.04u w=0.12u
m6286 VSS 4062 3272 VSS nch l=0.04u w=0.4u
m6287 3288 2508 3273 VSS nch l=0.04u w=0.4u
m6288 71211 3412 2909 VSS nch l=0.04u w=0.8u
m6289 3274 3336 71193 VSS nch l=0.04u w=0.8u
m6290 71212 3414 2911 VSS nch l=0.04u w=0.8u
m6291 3275 3337 71194 VSS nch l=0.04u w=0.8u
m6292 3276 3481 71195 VSS nch l=0.04u w=0.8u
m6293 3277 3482 71196 VSS nch l=0.04u w=0.8u
m6294 71213 3416 2913 VSS nch l=0.04u w=0.8u
m6295 3278 3338 71197 VSS nch l=0.04u w=0.8u
m6296 3279 131 71198 VSS nch l=0.04u w=0.8u
m6297 3280 3339 71199 VSS nch l=0.04u w=0.8u
m6298 71214 3420 2917 VSS nch l=0.04u w=0.8u
m6299 3281 3340 71200 VSS nch l=0.04u w=0.8u
m6300 3282 3341 71201 VSS nch l=0.04u w=0.8u
m6301 3283 3342 71202 VSS nch l=0.04u w=0.8u
m6302 71215 3424 2921 VSS nch l=0.04u w=0.8u
m6303 3284 3343 71203 VSS nch l=0.04u w=0.8u
m6304 3285 FBDIV[10] 71204 VSS nch l=0.04u w=0.8u
m6305 71216 3248 VSS VSS nch l=0.04u w=0.8u
m6306 3286 FBDIV[11] 71205 VSS nch l=0.04u w=0.8u
m6307 3291 4251 VSS VSS nch l=0.04u w=0.4u
m6308 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6309 VSS 3297 71206 VSS nch l=0.04u w=0.12u
m6310 VSS 3298 71207 VSS nch l=0.04u w=0.12u
m6311 VSS 3299 71208 VSS nch l=0.04u w=0.12u
m6312 VSS 3300 71209 VSS nch l=0.04u w=0.12u
m6313 2508 3273 3288 VSS nch l=0.04u w=0.4u
m6314 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6315 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6316 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6317 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6318 3293 3255 VSS VSS nch l=0.04u w=0.4u
m6319 3294 731 VSS VSS nch l=0.04u w=0.4u
m6320 VSS 3320 71211 VSS nch l=0.04u w=0.8u
m6321 VSS 3322 71212 VSS nch l=0.04u w=0.8u
m6322 VSS 3324 71213 VSS nch l=0.04u w=0.8u
m6323 VSS 3329 71214 VSS nch l=0.04u w=0.8u
m6324 VSS 3333 71215 VSS nch l=0.04u w=0.8u
m6325 3289 3198 71216 VSS nch l=0.04u w=0.8u
m6326 3295 4328 VSS VSS nch l=0.04u w=0.4u
m6327 71219 1676 3290 VSS nch l=0.04u w=0.8u
m6328 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6329 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6330 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6331 VSS 3287 3292 VSS nch l=0.04u w=0.4u
m6332 3296 4328 VSS VSS nch l=0.04u w=0.4u
m6333 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6334 3297 3266 VSS VSS nch l=0.04u w=0.4u
m6335 3298 3267 VSS VSS nch l=0.04u w=0.4u
m6336 3299 3268 VSS VSS nch l=0.04u w=0.4u
m6337 3300 3269 VSS VSS nch l=0.04u w=0.4u
m6338 3301 3318 2926 VSS nch l=0.04u w=0.4u
m6339 3302 110 3294 VSS nch l=0.04u w=0.4u
m6340 71220 3198 3289 VSS nch l=0.04u w=0.8u
m6341 3303 3336 VSS VSS nch l=0.04u w=0.4u
m6342 3304 3337 VSS VSS nch l=0.04u w=0.4u
m6343 3305 3276 VSS VSS nch l=0.04u w=0.4u
m6344 3306 3277 VSS VSS nch l=0.04u w=0.4u
m6345 3307 3338 VSS VSS nch l=0.04u w=0.4u
m6346 3308 131 VSS VSS nch l=0.04u w=0.4u
m6347 3309 3339 VSS VSS nch l=0.04u w=0.4u
m6348 3310 3340 VSS VSS nch l=0.04u w=0.4u
m6349 3311 3341 VSS VSS nch l=0.04u w=0.4u
m6350 3312 3342 VSS VSS nch l=0.04u w=0.4u
m6351 3313 3343 VSS VSS nch l=0.04u w=0.4u
m6352 3314 FBDIV[10] VSS VSS nch l=0.04u w=0.4u
m6353 VSS 4062 71219 VSS nch l=0.04u w=0.8u
m6354 71222 3250 VSS VSS nch l=0.04u w=0.8u
m6355 3316 3291 3212 VSS nch l=0.04u w=0.4u
m6356 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6357 415 3292 VSS VSS nch l=0.04u w=0.4u
m6358 3318 2926 3301 VSS nch l=0.04u w=0.4u
m6359 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6360 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6361 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6362 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6363 110 3294 3302 VSS nch l=0.04u w=0.4u
m6364 VSS 3248 71220 VSS nch l=0.04u w=0.8u
m6365 71223 3183 VSS VSS nch l=0.04u w=0.8u
m6366 3321 3338 3303 VSS nch l=0.04u w=0.4u
m6367 71224 3185 VSS VSS nch l=0.04u w=0.8u
m6368 3323 1908 3304 VSS nch l=0.04u w=0.4u
m6369 71225 3187 VSS VSS nch l=0.04u w=0.8u
m6370 3325 FRAC[10] 3307 VSS nch l=0.04u w=0.4u
m6371 3327 3339 3308 VSS nch l=0.04u w=0.4u
m6372 3328 3352 3309 VSS nch l=0.04u w=0.4u
m6373 71226 3191 VSS VSS nch l=0.04u w=0.8u
m6374 3330 3254 3310 VSS nch l=0.04u w=0.4u
m6375 3331 3265 3311 VSS nch l=0.04u w=0.4u
m6376 3332 3353 3312 VSS nch l=0.04u w=0.4u
m6377 71227 3195 VSS VSS nch l=0.04u w=0.8u
m6378 3334 FRAC[10] 3313 VSS nch l=0.04u w=0.4u
m6379 3335 3265 3314 VSS nch l=0.04u w=0.4u
m6380 3326 3295 3315 VSS nch l=0.04u w=0.4u
m6381 3317 3177 71222 VSS nch l=0.04u w=0.8u
m6382 71228 4251 3316 VSS nch l=0.04u w=0.12u
m6383 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6384 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6385 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6386 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6387 3345 3296 3234 VSS nch l=0.04u w=0.4u
m6388 3346 4328 3297 VSS nch l=0.04u w=0.4u
m6389 3347 4328 3298 VSS nch l=0.04u w=0.4u
m6390 3348 4328 3299 VSS nch l=0.04u w=0.4u
m6391 3349 4328 3300 VSS nch l=0.04u w=0.4u
m6392 71229 3288 3319 VSS nch l=0.04u w=0.8u
m6393 3320 3228 71223 VSS nch l=0.04u w=0.8u
m6394 3338 3303 3321 VSS nch l=0.04u w=0.4u
m6395 3322 3229 71224 VSS nch l=0.04u w=0.8u
m6396 1908 3304 3323 VSS nch l=0.04u w=0.4u
m6397 3324 3230 71225 VSS nch l=0.04u w=0.8u
m6398 FRAC[10] 3307 3325 VSS nch l=0.04u w=0.4u
m6399 3339 3308 3327 VSS nch l=0.04u w=0.4u
m6400 3352 3309 3328 VSS nch l=0.04u w=0.4u
m6401 3329 3231 71226 VSS nch l=0.04u w=0.8u
m6402 3254 3310 3330 VSS nch l=0.04u w=0.4u
m6403 3265 3311 3331 VSS nch l=0.04u w=0.4u
m6404 3353 3312 3332 VSS nch l=0.04u w=0.4u
m6405 3333 3232 71227 VSS nch l=0.04u w=0.8u
m6406 FRAC[10] 3313 3334 VSS nch l=0.04u w=0.4u
m6407 3265 3314 3335 VSS nch l=0.04u w=0.4u
m6408 3354 4328 VSS VSS nch l=0.04u w=0.4u
m6409 3355 4328 VSS VSS nch l=0.04u w=0.4u
m6410 3356 4328 VSS VSS nch l=0.04u w=0.4u
m6411 3357 4328 VSS VSS nch l=0.04u w=0.4u
m6412 71230 4328 3326 VSS nch l=0.04u w=0.12u
m6413 VSS 4062 3344 VSS nch l=0.04u w=0.4u
m6414 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6415 VSS 3364 71228 VSS nch l=0.04u w=0.12u
m6416 3358 4328 VSS VSS nch l=0.04u w=0.4u
m6417 71233 4328 3345 VSS nch l=0.04u w=0.12u
m6418 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6419 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6420 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6421 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6422 71234 3235 3346 VSS nch l=0.04u w=0.12u
m6423 71235 3236 3347 VSS nch l=0.04u w=0.12u
m6424 71236 3237 3348 VSS nch l=0.04u w=0.12u
m6425 71237 3238 3349 VSS nch l=0.04u w=0.12u
m6426 VSS 3318 3350 VSS nch l=0.04u w=0.4u
m6427 VSS 3115 71229 VSS nch l=0.04u w=0.8u
m6428 3359 4251 VSS VSS nch l=0.04u w=0.4u
m6429 VSS 3370 71230 VSS nch l=0.04u w=0.12u
m6430 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6431 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6432 3364 3316 VSS VSS nch l=0.04u w=0.4u
m6433 71254 3317 VSS VSS nch l=0.04u w=0.8u
m6434 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6435 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6436 VSS 3383 71233 VSS nch l=0.04u w=0.12u
m6437 VSS 3340 71234 VSS nch l=0.04u w=0.12u
m6438 VSS 3066 71235 VSS nch l=0.04u w=0.12u
m6439 VSS 3343 71236 VSS nch l=0.04u w=0.12u
m6440 VSS 3068 71237 VSS nch l=0.04u w=0.12u
m6441 71255 3302 3360 VSS nch l=0.04u w=0.8u
m6442 3370 3326 VSS VSS nch l=0.04u w=0.4u
m6443 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6444 3366 3354 3362 VSS nch l=0.04u w=0.4u
m6445 3367 3355 3363 VSS nch l=0.04u w=0.4u
m6446 3368 3356 3305 VSS nch l=0.04u w=0.4u
m6447 3369 3357 3306 VSS nch l=0.04u w=0.4u
m6448 3381 3386 3013 VSS nch l=0.04u w=0.4u
m6449 3365 3286 71254 VSS nch l=0.04u w=0.8u
m6450 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6451 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6452 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6453 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6454 3383 3345 VSS VSS nch l=0.04u w=0.4u
m6455 3382 3358 3287 VSS nch l=0.04u w=0.4u
m6456 3340 3346 VSS VSS nch l=0.04u w=0.4u
m6457 3066 3347 VSS VSS nch l=0.04u w=0.4u
m6458 3343 3348 VSS VSS nch l=0.04u w=0.4u
m6459 3068 3349 VSS VSS nch l=0.04u w=0.4u
m6460 71256 3953 3318 VSS nch l=0.04u w=0.8u
m6461 71257 3319 VSS VSS nch l=0.04u w=0.8u
m6462 VSS 3136 71255 VSS nch l=0.04u w=0.8u
m6463 3384 3359 3289 VSS nch l=0.04u w=0.4u
m6464 71259 4328 3366 VSS nch l=0.04u w=0.12u
m6465 71260 4328 3367 VSS nch l=0.04u w=0.12u
m6466 3228 3389 3204 VSS nch l=0.04u w=0.4u
m6467 71261 3321 3371 VSS nch l=0.04u w=0.8u
m6468 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6469 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6470 3229 3390 2024 VSS nch l=0.04u w=0.4u
m6471 71262 3323 3372 VSS nch l=0.04u w=0.8u
m6472 71263 4328 3368 VSS nch l=0.04u w=0.12u
m6473 71264 4328 3369 VSS nch l=0.04u w=0.12u
m6474 3230 3391 FRAC[14] VSS nch l=0.04u w=0.4u
m6475 71265 3325 3373 VSS nch l=0.04u w=0.8u
m6476 71266 3327 3374 VSS nch l=0.04u w=0.8u
m6477 71267 3328 3375 VSS nch l=0.04u w=0.8u
m6478 3231 3392 2744 VSS nch l=0.04u w=0.4u
m6479 71268 3330 3376 VSS nch l=0.04u w=0.8u
m6480 71269 3331 3377 VSS nch l=0.04u w=0.8u
m6481 71270 3332 3378 VSS nch l=0.04u w=0.8u
m6482 3232 3393 FRAC[14] VSS nch l=0.04u w=0.4u
m6483 71271 3334 3379 VSS nch l=0.04u w=0.8u
m6484 71272 3335 3380 VSS nch l=0.04u w=0.8u
m6485 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6486 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6487 3386 3013 3381 VSS nch l=0.04u w=0.4u
m6488 71273 3286 3365 VSS nch l=0.04u w=0.8u
m6489 3387 4251 3364 VSS nch l=0.04u w=0.4u
m6490 71274 4328 3382 VSS nch l=0.04u w=0.12u
m6491 VSS 3400 71256 VSS nch l=0.04u w=0.8u
m6492 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6493 3385 3227 71257 VSS nch l=0.04u w=0.8u
m6494 71276 4251 3384 VSS nch l=0.04u w=0.12u
m6495 VSS 3402 71259 VSS nch l=0.04u w=0.12u
m6496 VSS 3403 71260 VSS nch l=0.04u w=0.12u
m6497 3389 3204 3228 VSS nch l=0.04u w=0.4u
m6498 VSS 3145 71261 VSS nch l=0.04u w=0.8u
m6499 3390 2024 3229 VSS nch l=0.04u w=0.4u
m6500 VSS 3147 71262 VSS nch l=0.04u w=0.8u
m6501 VSS 3404 71263 VSS nch l=0.04u w=0.12u
m6502 VSS 3405 71264 VSS nch l=0.04u w=0.12u
m6503 3391 FRAC[14] 3230 VSS nch l=0.04u w=0.4u
m6504 VSS 3149 71265 VSS nch l=0.04u w=0.8u
m6505 3388 4328 3370 VSS nch l=0.04u w=0.4u
m6506 VSS 3150 71266 VSS nch l=0.04u w=0.8u
m6507 VSS 3151 71267 VSS nch l=0.04u w=0.8u
m6508 3392 2744 3231 VSS nch l=0.04u w=0.4u
m6509 VSS 3153 71268 VSS nch l=0.04u w=0.8u
m6510 VSS 3154 71269 VSS nch l=0.04u w=0.8u
m6511 VSS 3155 71270 VSS nch l=0.04u w=0.8u
m6512 3393 FRAC[14] 3232 VSS nch l=0.04u w=0.4u
m6513 VSS 3157 71271 VSS nch l=0.04u w=0.8u
m6514 VSS 3158 71272 VSS nch l=0.04u w=0.8u
m6515 VSS 3317 71273 VSS nch l=0.04u w=0.8u
m6516 71277 3291 3387 VSS nch l=0.04u w=0.12u
m6517 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6518 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6519 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6520 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6521 VSS 3406 71274 VSS nch l=0.04u w=0.12u
m6522 3395 4328 3383 VSS nch l=0.04u w=0.4u
m6523 3396 4328 VSS VSS nch l=0.04u w=0.4u
m6524 3397 4328 VSS VSS nch l=0.04u w=0.4u
m6525 3398 4328 VSS VSS nch l=0.04u w=0.4u
m6526 3399 4328 VSS VSS nch l=0.04u w=0.4u
m6527 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6528 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6529 VSS 3410 71276 VSS nch l=0.04u w=0.12u
m6530 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6531 71279 3360 VSS VSS nch l=0.04u w=0.8u
m6532 3402 3366 VSS VSS nch l=0.04u w=0.4u
m6533 3403 3367 VSS VSS nch l=0.04u w=0.4u
m6534 VSS 3203 3389 VSS nch l=0.04u w=0.4u
m6535 VSS 3208 3390 VSS nch l=0.04u w=0.4u
m6536 3404 3368 VSS VSS nch l=0.04u w=0.4u
m6537 3405 3369 VSS VSS nch l=0.04u w=0.4u
m6538 VSS 3204 3391 VSS nch l=0.04u w=0.4u
m6539 71280 3295 3388 VSS nch l=0.04u w=0.12u
m6540 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6541 VSS 2854 3392 VSS nch l=0.04u w=0.4u
m6542 VSS 2856 3393 VSS nch l=0.04u w=0.4u
m6543 VSS 3386 3394 VSS nch l=0.04u w=0.4u
m6544 VSS 3070 71277 VSS nch l=0.04u w=0.12u
m6545 3406 3382 VSS VSS nch l=0.04u w=0.4u
m6546 71281 3296 3395 VSS nch l=0.04u w=0.12u
m6547 VSS 3434 3400 VSS nch l=0.04u w=0.4u
m6548 VSS 3179 VSS VSS nch l=0.26u w=0.8u
m6549 3410 3384 VSS VSS nch l=0.04u w=0.4u
m6550 3411 3288 VSS VSS nch l=0.04u w=0.4u
m6551 3401 3256 71279 VSS nch l=0.04u w=0.8u
m6552 VSS 3440 71280 VSS nch l=0.04u w=0.12u
m6553 71282 3371 VSS VSS nch l=0.04u w=0.8u
m6554 71283 3372 VSS VSS nch l=0.04u w=0.8u
m6555 71284 3373 VSS VSS nch l=0.04u w=0.8u
m6556 71285 3374 VSS VSS nch l=0.04u w=0.8u
m6557 71286 3375 VSS VSS nch l=0.04u w=0.8u
m6558 71287 3376 VSS VSS nch l=0.04u w=0.8u
m6559 71288 3377 VSS VSS nch l=0.04u w=0.8u
m6560 71289 3378 VSS VSS nch l=0.04u w=0.8u
m6561 71290 3379 VSS VSS nch l=0.04u w=0.8u
m6562 71291 3380 VSS VSS nch l=0.04u w=0.8u
m6563 3070 3387 VSS VSS nch l=0.04u w=0.4u
m6564 3427 4251 VSS VSS nch l=0.04u w=0.4u
m6565 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6566 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6567 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6568 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6569 VSS 3442 71281 VSS nch l=0.04u w=0.12u
m6570 3428 3396 3407 VSS nch l=0.04u w=0.4u
m6571 3429 3397 3408 VSS nch l=0.04u w=0.4u
m6572 3430 3398 3409 VSS nch l=0.04u w=0.4u
m6573 3431 3399 3341 VSS nch l=0.04u w=0.4u
m6574 3432 3433 VSS VSS nch l=0.04u w=0.8u
m6575 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6576 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6577 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6578 VSS 3209 VSS VSS nch l=0.26u w=0.8u
m6579 3435 3115 3411 VSS nch l=0.04u w=0.4u
m6580 3440 3388 VSS VSS nch l=0.04u w=0.4u
m6581 3436 4328 3402 VSS nch l=0.04u w=0.4u
m6582 3437 4328 3403 VSS nch l=0.04u w=0.4u
m6583 71293 3203 3412 VSS nch l=0.04u w=0.8u
m6584 3413 3274 71282 VSS nch l=0.04u w=0.8u
m6585 71294 3208 3414 VSS nch l=0.04u w=0.8u
m6586 3415 3275 71283 VSS nch l=0.04u w=0.8u
m6587 3438 4328 3404 VSS nch l=0.04u w=0.4u
m6588 3439 4328 3405 VSS nch l=0.04u w=0.4u
m6589 71295 3204 3416 VSS nch l=0.04u w=0.8u
m6590 3417 3278 71284 VSS nch l=0.04u w=0.8u
m6591 3418 3279 71285 VSS nch l=0.04u w=0.8u
m6592 3419 3280 71286 VSS nch l=0.04u w=0.8u
m6593 71296 2854 3420 VSS nch l=0.04u w=0.8u
m6594 3421 3281 71287 VSS nch l=0.04u w=0.8u
m6595 3422 3282 71288 VSS nch l=0.04u w=0.8u
m6596 3423 3283 71289 VSS nch l=0.04u w=0.8u
m6597 71297 2856 3424 VSS nch l=0.04u w=0.8u
m6598 3425 3284 71290 VSS nch l=0.04u w=0.8u
m6599 3426 3285 71291 VSS nch l=0.04u w=0.8u
m6600 71298 3953 3386 VSS nch l=0.04u w=0.8u
m6601 3442 3395 VSS VSS nch l=0.04u w=0.4u
m6602 3441 4328 3406 VSS nch l=0.04u w=0.4u
m6603 71299 4328 3428 VSS nch l=0.04u w=0.12u
m6604 71300 4328 3429 VSS nch l=0.04u w=0.12u
m6605 71301 4328 3430 VSS nch l=0.04u w=0.12u
m6606 71302 4328 3431 VSS nch l=0.04u w=0.12u
m6607 71303 3484 3434 VSS nch l=0.04u w=0.8u
m6608 3446 3445 VSS VSS nch l=0.04u w=0.8u
m6609 3115 3411 3435 VSS nch l=0.04u w=0.4u
m6610 3447 4251 3410 VSS nch l=0.04u w=0.4u
m6611 3448 3302 VSS VSS nch l=0.04u w=0.4u
m6612 71304 3354 3436 VSS nch l=0.04u w=0.12u
m6613 71305 3355 3437 VSS nch l=0.04u w=0.12u
m6614 VSS 3204 71293 VSS nch l=0.04u w=0.8u
m6615 VSS 2024 71294 VSS nch l=0.04u w=0.8u
m6616 71306 3356 3438 VSS nch l=0.04u w=0.12u
m6617 71307 3357 3439 VSS nch l=0.04u w=0.12u
m6618 VSS FRAC[14] 71295 VSS nch l=0.04u w=0.8u
m6619 VSS 2744 71296 VSS nch l=0.04u w=0.8u
m6620 VSS FRAC[14] 71297 VSS nch l=0.04u w=0.8u
m6621 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6622 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6623 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6624 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6625 VSS 3484 71298 VSS nch l=0.04u w=0.8u
m6626 3450 3070 VSS VSS nch l=0.04u w=0.4u
m6627 3449 3427 3365 VSS nch l=0.04u w=0.4u
m6628 71309 3358 3441 VSS nch l=0.04u w=0.12u
m6629 VSS 3470 71299 VSS nch l=0.04u w=0.12u
m6630 VSS 3471 71300 VSS nch l=0.04u w=0.12u
m6631 VSS 3472 71301 VSS nch l=0.04u w=0.12u
m6632 VSS 3473 71302 VSS nch l=0.04u w=0.12u
m6633 VSS 3240 VSS VSS nch l=0.26u w=0.8u
m6634 VSS 3241 VSS VSS nch l=0.26u w=0.8u
m6635 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6636 71310 4351 71303 VSS nch l=0.04u w=0.8u
m6637 VSS 3443 3443 VSS nch l=0.04u w=0.8u
m6638 71311 3359 3447 VSS nch l=0.04u w=0.12u
m6639 3454 3136 3448 VSS nch l=0.04u w=0.4u
m6640 VSS 3478 71304 VSS nch l=0.04u w=0.12u
m6641 VSS 3336 71305 VSS nch l=0.04u w=0.12u
m6642 VSS 3479 71306 VSS nch l=0.04u w=0.12u
m6643 VSS 3338 71307 VSS nch l=0.04u w=0.12u
m6644 3456 3321 VSS VSS nch l=0.04u w=0.4u
m6645 3458 3323 VSS VSS nch l=0.04u w=0.4u
m6646 3460 3325 VSS VSS nch l=0.04u w=0.4u
m6647 3461 3327 VSS VSS nch l=0.04u w=0.4u
m6648 3462 3328 VSS VSS nch l=0.04u w=0.4u
m6649 3464 3330 VSS VSS nch l=0.04u w=0.4u
m6650 3465 3331 VSS VSS nch l=0.04u w=0.4u
m6651 3466 3332 VSS VSS nch l=0.04u w=0.4u
m6652 3468 3334 VSS VSS nch l=0.04u w=0.4u
m6653 3469 3335 VSS VSS nch l=0.04u w=0.4u
m6654 VSS 3070 3450 VSS nch l=0.04u w=0.4u
m6655 71314 4251 3449 VSS nch l=0.04u w=0.12u
m6656 VSS 3485 71309 VSS nch l=0.04u w=0.12u
m6657 VSS 3442 3451 VSS nch l=0.04u w=0.4u
m6658 3470 3428 VSS VSS nch l=0.04u w=0.4u
m6659 3471 3429 VSS VSS nch l=0.04u w=0.4u
m6660 3472 3430 VSS VSS nch l=0.04u w=0.4u
m6661 3473 3431 VSS VSS nch l=0.04u w=0.4u
m6662 3474 3475 VSS VSS nch l=0.04u w=0.8u
m6663 3477 3476 VSS VSS nch l=0.04u w=0.8u
m6664 VSS 3490 71310 VSS nch l=0.04u w=0.8u
m6665 VSS 3453 3453 VSS nch l=0.04u w=0.8u
m6666 VSS 3122 71311 VSS nch l=0.04u w=0.12u
m6667 3136 3448 3454 VSS nch l=0.04u w=0.4u
m6668 3478 3436 VSS VSS nch l=0.04u w=0.4u
m6669 3336 3437 VSS VSS nch l=0.04u w=0.4u
m6670 VSS 3258 VSS VSS nch l=0.26u w=0.8u
m6671 VSS 3259 VSS VSS nch l=0.26u w=0.8u
m6672 3479 3438 VSS VSS nch l=0.04u w=0.4u
m6673 3338 3439 VSS VSS nch l=0.04u w=0.4u
m6674 VSS 3262 VSS VSS nch l=0.26u w=0.8u
m6675 VSS 3263 VSS VSS nch l=0.26u w=0.8u
m6676 3480 2445 VSS VSS nch l=0.04u w=0.4u
m6677 3363 3145 3456 VSS nch l=0.04u w=0.4u
m6678 3482 3147 3458 VSS nch l=0.04u w=0.4u
m6679 3337 3149 3460 VSS nch l=0.04u w=0.4u
m6680 3315 3150 3461 VSS nch l=0.04u w=0.4u
m6681 3408 3151 3462 VSS nch l=0.04u w=0.4u
m6682 3253 3153 3464 VSS nch l=0.04u w=0.4u
m6683 3352 3154 3465 VSS nch l=0.04u w=0.4u
m6684 3341 3155 3466 VSS nch l=0.04u w=0.4u
m6685 3254 3157 3468 VSS nch l=0.04u w=0.4u
m6686 3353 3158 3469 VSS nch l=0.04u w=0.4u
m6687 VSS 3505 71314 VSS nch l=0.04u w=0.12u
m6688 3484 3518 VSS VSS nch l=0.04u w=0.4u
m6689 3485 3441 VSS VSS nch l=0.04u w=0.4u
m6690 1321 3451 VSS VSS nch l=0.04u w=0.4u
m6691 VSS 3270 VSS VSS nch l=0.26u w=0.8u
m6692 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m6693 3122 3447 VSS VSS nch l=0.04u w=0.4u
m6694 3491 3492 VSS VSS nch l=0.04u w=0.8u
m6695 3494 3493 VSS VSS nch l=0.04u w=0.8u
m6696 3495 3496 VSS VSS nch l=0.04u w=0.8u
m6697 3498 3497 VSS VSS nch l=0.04u w=0.8u
m6698 VSS 3435 3480 VSS nch l=0.04u w=0.4u
m6699 3499 3385 VSS VSS nch l=0.04u w=0.4u
m6700 3145 3456 3363 VSS nch l=0.04u w=0.4u
m6701 3147 3458 3482 VSS nch l=0.04u w=0.4u
m6702 3149 3460 3337 VSS nch l=0.04u w=0.4u
m6703 3150 3461 3315 VSS nch l=0.04u w=0.4u
m6704 3151 3462 3408 VSS nch l=0.04u w=0.4u
m6705 3153 3464 3253 VSS nch l=0.04u w=0.4u
m6706 3154 3465 3352 VSS nch l=0.04u w=0.4u
m6707 3155 3466 3341 VSS nch l=0.04u w=0.4u
m6708 3157 3468 3254 VSS nch l=0.04u w=0.4u
m6709 3158 3469 3353 VSS nch l=0.04u w=0.4u
m6710 3362 3513 3455 VSS nch l=0.04u w=0.4u
m6711 3481 3514 3457 VSS nch l=0.04u w=0.4u
m6712 3483 3515 3459 VSS nch l=0.04u w=0.4u
m6713 3086 3516 3463 VSS nch l=0.04u w=0.4u
m6714 3087 3517 3467 VSS nch l=0.04u w=0.4u
m6715 3505 3449 VSS VSS nch l=0.04u w=0.4u
m6716 VSS 3518 3484 VSS nch l=0.04u w=0.4u
m6717 71327 3450 VSS VSS nch l=0.04u w=0.8u
m6718 3512 3511 VSS VSS nch l=0.04u w=0.8u
m6719 3507 4328 3470 VSS nch l=0.04u w=0.4u
m6720 3508 4328 3471 VSS nch l=0.04u w=0.4u
m6721 3509 4328 3472 VSS nch l=0.04u w=0.4u
m6722 3510 4328 3473 VSS nch l=0.04u w=0.4u
m6723 VSS 3486 3486 VSS nch l=0.04u w=0.8u
m6724 VSS 3489 3489 VSS nch l=0.04u w=0.8u
m6725 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m6726 VSS 3523 3490 VSS nch l=0.04u w=0.4u
m6727 3513 3455 3362 VSS nch l=0.04u w=0.4u
m6728 3514 3457 3481 VSS nch l=0.04u w=0.4u
m6729 3515 3459 3483 VSS nch l=0.04u w=0.4u
m6730 3516 3463 3086 VSS nch l=0.04u w=0.4u
m6731 3517 3467 3087 VSS nch l=0.04u w=0.4u
m6732 71329 2969 71327 VSS nch l=0.04u w=0.8u
m6733 3519 4328 VSS VSS nch l=0.04u w=0.4u
m6734 3520 4328 VSS VSS nch l=0.04u w=0.4u
m6735 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m6736 71347 3396 3507 VSS nch l=0.04u w=0.12u
m6737 71348 3397 3508 VSS nch l=0.04u w=0.12u
m6738 71349 3398 3509 VSS nch l=0.04u w=0.12u
m6739 71350 3399 3510 VSS nch l=0.04u w=0.12u
m6740 3524 3122 VSS VSS nch l=0.04u w=0.4u
m6741 71353 2491 VSS VSS nch l=0.04u w=0.8u
m6742 71354 110 VSS VSS nch l=0.04u w=0.8u
m6743 VSS 3500 3513 VSS nch l=0.04u w=0.4u
m6744 VSS 3501 3514 VSS nch l=0.04u w=0.4u
m6745 VSS 3502 3515 VSS nch l=0.04u w=0.4u
m6746 VSS 3503 3516 VSS nch l=0.04u w=0.4u
m6747 VSS 3504 3517 VSS nch l=0.04u w=0.4u
m6748 3506 3484 71329 VSS nch l=0.04u w=0.8u
m6749 3527 4251 3505 VSS nch l=0.04u w=0.4u
m6750 VSS 3556 3518 VSS nch l=0.04u w=0.4u
m6751 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m6752 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m6753 VSS 3553 71347 VSS nch l=0.04u w=0.12u
m6754 VSS 3339 71348 VSS nch l=0.04u w=0.12u
m6755 VSS 3554 71349 VSS nch l=0.04u w=0.12u
m6756 VSS 3342 71350 VSS nch l=0.04u w=0.12u
m6757 VSS 3522 3522 VSS nch l=0.04u w=0.8u
m6758 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m6759 71355 4064 3523 VSS nch l=0.04u w=0.8u
m6760 VSS 3122 3524 VSS nch l=0.04u w=0.4u
m6761 71358 2739 71353 VSS nch l=0.04u w=0.8u
m6762 3526 1023 71354 VSS nch l=0.04u w=0.8u
m6763 VSS 3528 3528 VSS nch l=0.04u w=0.8u
m6764 VSS 3531 3531 VSS nch l=0.04u w=0.8u
m6765 71359 3610 VSS VSS nch l=0.04u w=0.8u
m6766 71360 1935 VSS VSS nch l=0.04u w=0.8u
m6767 71361 2616 VSS VSS nch l=0.04u w=0.8u
m6768 71362 2616 VSS VSS nch l=0.04u w=0.8u
m6769 VSS 3532 3532 VSS nch l=0.04u w=0.8u
m6770 VSS 3535 3535 VSS nch l=0.04u w=0.8u
m6771 71363 FRAC[11] VSS VSS nch l=0.04u w=0.8u
m6772 VSS 3582 3536 VSS nch l=0.04u w=0.4u
m6773 71364 3611 VSS VSS nch l=0.04u w=0.8u
m6774 71365 3622 VSS VSS nch l=0.04u w=0.8u
m6775 71366 3588 VSS VSS nch l=0.04u w=0.8u
m6776 71367 3536 VSS VSS nch l=0.04u w=0.8u
m6777 71368 3623 VSS VSS nch l=0.04u w=0.8u
m6778 71369 FRAC[11] VSS VSS nch l=0.04u w=0.8u
m6779 71370 3536 VSS VSS nch l=0.04u w=0.8u
m6780 71371 3427 3527 VSS nch l=0.04u w=0.12u
m6781 71372 3518 VSS VSS nch l=0.04u w=0.12u
m6782 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m6783 VSS 3538 3538 VSS nch l=0.04u w=0.8u
m6784 3551 3519 3485 VSS nch l=0.04u w=0.4u
m6785 3552 3520 3442 VSS nch l=0.04u w=0.4u
m6786 3553 3507 VSS VSS nch l=0.04u w=0.4u
m6787 3339 3508 VSS VSS nch l=0.04u w=0.4u
m6788 3554 3509 VSS VSS nch l=0.04u w=0.4u
m6789 3342 3510 VSS VSS nch l=0.04u w=0.4u
m6790 VSS 3565 71355 VSS nch l=0.04u w=0.8u
m6791 3525 3016 71358 VSS nch l=0.04u w=0.8u
m6792 71374 3693 3183 VSS nch l=0.04u w=0.8u
m6793 3539 3608 71359 VSS nch l=0.04u w=0.8u
m6794 71375 3695 3185 VSS nch l=0.04u w=0.8u
m6795 3540 3609 71360 VSS nch l=0.04u w=0.8u
m6796 3541 3761 71361 VSS nch l=0.04u w=0.8u
m6797 3542 3762 71362 VSS nch l=0.04u w=0.8u
m6798 71376 3697 3187 VSS nch l=0.04u w=0.8u
m6799 3543 3610 71363 VSS nch l=0.04u w=0.8u
m6800 3544 131 71364 VSS nch l=0.04u w=0.8u
m6801 3545 3611 71365 VSS nch l=0.04u w=0.8u
m6802 71377 3701 3191 VSS nch l=0.04u w=0.8u
m6803 3546 3612 71366 VSS nch l=0.04u w=0.8u
m6804 3547 3589 71367 VSS nch l=0.04u w=0.8u
m6805 3548 3613 71368 VSS nch l=0.04u w=0.8u
m6806 71378 3705 3195 VSS nch l=0.04u w=0.8u
m6807 3549 3614 71369 VSS nch l=0.04u w=0.8u
m6808 3550 FBDIV[11] 71370 VSS nch l=0.04u w=0.8u
m6809 VSS 3199 71371 VSS nch l=0.04u w=0.12u
m6810 3556 3660 71372 VSS nch l=0.04u w=0.12u
m6811 3555 3506 VSS VSS nch l=0.04u w=0.4u
m6812 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m6813 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m6814 VSS 3521 VSS VSS nch l=0.26u w=0.8u
m6815 71379 4328 3551 VSS nch l=0.04u w=0.12u
m6816 71380 4328 3552 VSS nch l=0.04u w=0.12u
m6817 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m6818 3557 3567 VSS VSS nch l=0.04u w=0.4u
m6819 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m6820 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m6821 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m6822 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m6823 3558 1023 VSS VSS nch l=0.04u w=0.4u
m6824 VSS 3591 71374 VSS nch l=0.04u w=0.8u
m6825 VSS 3593 71375 VSS nch l=0.04u w=0.8u
m6826 VSS 3595 71376 VSS nch l=0.04u w=0.8u
m6827 VSS 3600 71377 VSS nch l=0.04u w=0.8u
m6828 VSS 3604 71378 VSS nch l=0.04u w=0.8u
m6829 3199 3527 VSS VSS nch l=0.04u w=0.4u
m6830 3559 4328 VSS VSS nch l=0.04u w=0.4u
m6831 3560 4251 3556 VSS nch l=0.04u w=0.4u
m6832 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m6833 VSS 3537 VSS VSS nch l=0.26u w=0.8u
m6834 VSS 3584 71379 VSS nch l=0.04u w=0.12u
m6835 VSS 3585 71380 VSS nch l=0.04u w=0.12u
m6836 3561 4328 VSS VSS nch l=0.04u w=0.4u
m6837 3562 4328 VSS VSS nch l=0.04u w=0.4u
m6838 3563 4328 VSS VSS nch l=0.04u w=0.4u
m6839 3564 4328 VSS VSS nch l=0.04u w=0.4u
m6840 3565 3619 VSS VSS nch l=0.04u w=0.4u
m6841 3568 3525 VSS VSS nch l=0.04u w=0.4u
m6842 3569 110 3558 VSS nch l=0.04u w=0.4u
m6843 3570 3608 VSS VSS nch l=0.04u w=0.4u
m6844 3571 3609 VSS VSS nch l=0.04u w=0.4u
m6845 3572 3541 VSS VSS nch l=0.04u w=0.4u
m6846 3573 3542 VSS VSS nch l=0.04u w=0.4u
m6847 3574 3610 VSS VSS nch l=0.04u w=0.4u
m6848 3575 131 VSS VSS nch l=0.04u w=0.4u
m6849 3576 3611 VSS VSS nch l=0.04u w=0.4u
m6850 3577 3612 VSS VSS nch l=0.04u w=0.4u
m6851 3578 3589 VSS VSS nch l=0.04u w=0.4u
m6852 3579 3613 VSS VSS nch l=0.04u w=0.4u
m6853 3580 3614 VSS VSS nch l=0.04u w=0.4u
m6854 3581 FBDIV[11] VSS VSS nch l=0.04u w=0.4u
m6855 71383 3555 VSS VSS nch l=0.04u w=0.8u
m6856 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m6857 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m6858 VSS 3521 VSS VSS nch l=0.26u w=0.8u
m6859 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m6860 3584 3551 VSS VSS nch l=0.04u w=0.4u
m6861 3585 3552 VSS VSS nch l=0.04u w=0.4u
m6862 VSS 3619 3565 VSS nch l=0.04u w=0.4u
m6863 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m6864 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m6865 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m6866 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m6867 3566 3590 3567 VSS nch l=0.04u w=0.4u
m6868 110 3558 3569 VSS nch l=0.04u w=0.4u
m6869 71384 3455 VSS VSS nch l=0.04u w=0.8u
m6870 3592 3610 3570 VSS nch l=0.04u w=0.4u
m6871 71385 3457 VSS VSS nch l=0.04u w=0.8u
m6872 3594 1935 3571 VSS nch l=0.04u w=0.4u
m6873 71386 3459 VSS VSS nch l=0.04u w=0.8u
m6874 3596 FRAC[11] 3574 VSS nch l=0.04u w=0.4u
m6875 3598 3611 3575 VSS nch l=0.04u w=0.4u
m6876 3599 3622 3576 VSS nch l=0.04u w=0.4u
m6877 71387 3463 VSS VSS nch l=0.04u w=0.8u
m6878 3601 3588 3577 VSS nch l=0.04u w=0.4u
m6879 3602 3536 3578 VSS nch l=0.04u w=0.4u
m6880 3603 3623 3579 VSS nch l=0.04u w=0.4u
m6881 71388 3467 VSS VSS nch l=0.04u w=0.8u
m6882 3605 FRAC[11] 3580 VSS nch l=0.04u w=0.4u
m6883 3606 3536 3581 VSS nch l=0.04u w=0.4u
m6884 3607 3199 VSS VSS nch l=0.04u w=0.4u
m6885 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m6886 VSS 3537 VSS VSS nch l=0.26u w=0.8u
m6887 3597 3559 3582 VSS nch l=0.04u w=0.4u
m6888 VSS 3634 3560 VSS nch l=0.04u w=0.4u
m6889 3583 3953 71383 VSS nch l=0.04u w=0.8u
m6890 3615 3561 3586 VSS nch l=0.04u w=0.4u
m6891 3616 3562 3587 VSS nch l=0.04u w=0.4u
m6892 3617 3563 3588 VSS nch l=0.04u w=0.4u
m6893 3618 3564 3589 VSS nch l=0.04u w=0.4u
m6894 3590 3567 3566 VSS nch l=0.04u w=0.4u
m6895 71389 3568 VSS VSS nch l=0.04u w=0.8u
m6896 3591 3500 71384 VSS nch l=0.04u w=0.8u
m6897 3610 3570 3592 VSS nch l=0.04u w=0.4u
m6898 3593 3501 71385 VSS nch l=0.04u w=0.8u
m6899 1935 3571 3594 VSS nch l=0.04u w=0.4u
m6900 3595 3502 71386 VSS nch l=0.04u w=0.8u
m6901 FRAC[11] 3574 3596 VSS nch l=0.04u w=0.4u
m6902 3611 3575 3598 VSS nch l=0.04u w=0.4u
m6903 3622 3576 3599 VSS nch l=0.04u w=0.4u
m6904 3600 3503 71387 VSS nch l=0.04u w=0.8u
m6905 3588 3577 3601 VSS nch l=0.04u w=0.4u
m6906 3536 3578 3602 VSS nch l=0.04u w=0.4u
m6907 3623 3579 3603 VSS nch l=0.04u w=0.4u
m6908 3604 3504 71388 VSS nch l=0.04u w=0.8u
m6909 FRAC[11] 3580 3605 VSS nch l=0.04u w=0.4u
m6910 3536 3581 3606 VSS nch l=0.04u w=0.4u
m6911 VSS 3199 3607 VSS nch l=0.04u w=0.4u
m6912 3624 4328 VSS VSS nch l=0.04u w=0.4u
m6913 3625 4328 VSS VSS nch l=0.04u w=0.4u
m6914 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m6915 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m6916 3626 4328 VSS VSS nch l=0.04u w=0.4u
m6917 3627 4328 VSS VSS nch l=0.04u w=0.4u
m6918 71390 4328 3597 VSS nch l=0.04u w=0.12u
m6919 71391 3560 VSS VSS nch l=0.04u w=0.12u
m6920 VSS 3521 VSS VSS nch l=0.26u w=0.8u
m6921 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m6922 3628 4328 3584 VSS nch l=0.04u w=0.4u
m6923 3629 4328 3585 VSS nch l=0.04u w=0.4u
m6924 71393 4328 3615 VSS nch l=0.04u w=0.12u
m6925 71394 4328 3616 VSS nch l=0.04u w=0.12u
m6926 71395 4328 3617 VSS nch l=0.04u w=0.12u
m6927 71396 4328 3618 VSS nch l=0.04u w=0.12u
m6928 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m6929 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m6930 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m6931 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m6932 VSS 3659 3619 VSS nch l=0.04u w=0.4u
m6933 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m6934 VSS 3537 VSS VSS nch l=0.26u w=0.8u
m6935 71397 3288 71389 VSS nch l=0.04u w=0.8u
m6936 VSS 3641 71390 VSS nch l=0.04u w=0.12u
m6937 3634 4251 71391 VSS nch l=0.04u w=0.12u
m6938 3635 3583 VSS VSS nch l=0.04u w=0.4u
m6939 71413 3519 3628 VSS nch l=0.04u w=0.12u
m6940 71414 3520 3629 VSS nch l=0.04u w=0.12u
m6941 VSS 3655 71393 VSS nch l=0.04u w=0.12u
m6942 VSS 3656 71394 VSS nch l=0.04u w=0.12u
m6943 VSS 3657 71395 VSS nch l=0.04u w=0.12u
m6944 VSS 3658 71396 VSS nch l=0.04u w=0.12u
m6945 71415 3619 VSS VSS nch l=0.04u w=0.12u
m6946 3636 4062 VSS VSS nch l=0.04u w=0.4u
m6947 3620 2630 71397 VSS nch l=0.04u w=0.8u
m6948 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m6949 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m6950 VSS 3521 VSS VSS nch l=0.26u w=0.8u
m6951 71416 3569 3630 VSS nch l=0.04u w=0.8u
m6952 3641 3597 VSS VSS nch l=0.04u w=0.4u
m6953 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m6954 3642 3660 3634 VSS nch l=0.04u w=0.4u
m6955 3643 3484 VSS VSS nch l=0.04u w=0.4u
m6956 3637 3624 3632 VSS nch l=0.04u w=0.4u
m6957 3638 3625 3633 VSS nch l=0.04u w=0.4u
m6958 3639 3626 3572 VSS nch l=0.04u w=0.4u
m6959 3640 3627 3573 VSS nch l=0.04u w=0.4u
m6960 VSS 3662 71413 VSS nch l=0.04u w=0.12u
m6961 VSS 3663 71414 VSS nch l=0.04u w=0.12u
m6962 3655 3615 VSS VSS nch l=0.04u w=0.4u
m6963 3656 3616 VSS VSS nch l=0.04u w=0.4u
m6964 3657 3617 VSS VSS nch l=0.04u w=0.4u
m6965 3658 3618 VSS VSS nch l=0.04u w=0.4u
m6966 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m6967 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m6968 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m6969 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m6970 3659 3756 71415 VSS nch l=0.04u w=0.12u
m6971 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m6972 VSS 3537 VSS VSS nch l=0.26u w=0.8u
m6973 VSS 3401 71416 VSS nch l=0.04u w=0.8u
m6974 71417 4328 3637 VSS nch l=0.04u w=0.12u
m6975 71418 4328 3638 VSS nch l=0.04u w=0.12u
m6976 3500 3668 3479 VSS nch l=0.04u w=0.4u
m6977 71419 3592 3644 VSS nch l=0.04u w=0.8u
m6978 3501 3669 1998 VSS nch l=0.04u w=0.4u
m6979 71420 3594 3645 VSS nch l=0.04u w=0.8u
m6980 71421 4328 3639 VSS nch l=0.04u w=0.12u
m6981 71422 4328 3640 VSS nch l=0.04u w=0.12u
m6982 3502 3670 FRAC[13] VSS nch l=0.04u w=0.4u
m6983 71423 3596 3646 VSS nch l=0.04u w=0.8u
m6984 71424 3598 3647 VSS nch l=0.04u w=0.8u
m6985 71425 3599 3648 VSS nch l=0.04u w=0.8u
m6986 3503 3671 3087 VSS nch l=0.04u w=0.4u
m6987 71426 3601 3649 VSS nch l=0.04u w=0.8u
m6988 71427 3602 3650 VSS nch l=0.04u w=0.8u
m6989 71428 3603 3651 VSS nch l=0.04u w=0.8u
m6990 3504 3672 FRAC[13] VSS nch l=0.04u w=0.4u
m6991 71429 3605 3652 VSS nch l=0.04u w=0.8u
m6992 71430 3606 3653 VSS nch l=0.04u w=0.8u
m6993 3654 3661 3583 VSS nch l=0.04u w=0.4u
m6994 3662 3628 VSS VSS nch l=0.04u w=0.4u
m6995 3663 3629 VSS VSS nch l=0.04u w=0.4u
m6996 3664 4251 3659 VSS nch l=0.04u w=0.4u
m6997 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m6998 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m6999 VSS 3521 VSS VSS nch l=0.26u w=0.8u
m7000 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m7001 71431 4062 VSS VSS nch l=0.04u w=0.8u
m7002 71432 3499 VSS VSS nch l=0.04u w=0.8u
m7003 VSS 3681 71417 VSS nch l=0.04u w=0.12u
m7004 VSS 3682 71418 VSS nch l=0.04u w=0.12u
m7005 3668 3479 3500 VSS nch l=0.04u w=0.4u
m7006 VSS 3413 71419 VSS nch l=0.04u w=0.8u
m7007 3669 1998 3501 VSS nch l=0.04u w=0.4u
m7008 VSS 3415 71420 VSS nch l=0.04u w=0.8u
m7009 VSS 3683 71421 VSS nch l=0.04u w=0.12u
m7010 VSS 3684 71422 VSS nch l=0.04u w=0.12u
m7011 3670 FRAC[13] 3502 VSS nch l=0.04u w=0.4u
m7012 VSS 3417 71423 VSS nch l=0.04u w=0.8u
m7013 3667 4328 3641 VSS nch l=0.04u w=0.4u
m7014 VSS 3418 71424 VSS nch l=0.04u w=0.8u
m7015 VSS 3419 71425 VSS nch l=0.04u w=0.8u
m7016 3671 3087 3503 VSS nch l=0.04u w=0.4u
m7017 VSS 3421 71426 VSS nch l=0.04u w=0.8u
m7018 VSS 3422 71427 VSS nch l=0.04u w=0.8u
m7019 VSS 3423 71428 VSS nch l=0.04u w=0.8u
m7020 3672 FRAC[13] 3504 VSS nch l=0.04u w=0.4u
m7021 VSS 3425 71429 VSS nch l=0.04u w=0.8u
m7022 VSS 3426 71430 VSS nch l=0.04u w=0.8u
m7023 VSS 4251 3660 VSS nch l=0.04u w=0.4u
m7024 71433 3607 VSS VSS nch l=0.04u w=0.8u
m7025 3661 3583 3654 VSS nch l=0.04u w=0.4u
m7026 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m7027 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m7028 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m7029 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m7030 3674 4328 3655 VSS nch l=0.04u w=0.4u
m7031 3675 4328 3656 VSS nch l=0.04u w=0.4u
m7032 3676 4328 3657 VSS nch l=0.04u w=0.4u
m7033 3677 4328 3658 VSS nch l=0.04u w=0.4u
m7034 VSS 3444 VSS VSS nch l=0.26u w=0.8u
m7035 VSS 3537 VSS VSS nch l=0.26u w=0.8u
m7036 3679 3678 VSS VSS nch l=0.04u w=0.8u
m7037 3665 616 71431 VSS nch l=0.04u w=0.8u
m7038 3666 3620 71432 VSS nch l=0.04u w=0.8u
m7039 71434 3630 VSS VSS nch l=0.04u w=0.8u
m7040 3681 3637 VSS VSS nch l=0.04u w=0.4u
m7041 3682 3638 VSS VSS nch l=0.04u w=0.4u
m7042 VSS 3478 3668 VSS nch l=0.04u w=0.4u
m7043 VSS 3483 3669 VSS nch l=0.04u w=0.4u
m7044 3683 3639 VSS VSS nch l=0.04u w=0.4u
m7045 3684 3640 VSS VSS nch l=0.04u w=0.4u
m7046 VSS 3479 3670 VSS nch l=0.04u w=0.4u
m7047 71435 3559 3667 VSS nch l=0.04u w=0.12u
m7048 VSS 3201 3671 VSS nch l=0.04u w=0.4u
m7049 VSS 3202 3672 VSS nch l=0.04u w=0.4u
m7050 71436 3017 71433 VSS nch l=0.04u w=0.8u
m7051 3685 4328 VSS VSS nch l=0.04u w=0.4u
m7052 3686 4328 VSS VSS nch l=0.04u w=0.4u
m7053 71437 3561 3674 VSS nch l=0.04u w=0.12u
m7054 71438 3562 3675 VSS nch l=0.04u w=0.12u
m7055 71439 3563 3676 VSS nch l=0.04u w=0.12u
m7056 71440 3564 3677 VSS nch l=0.04u w=0.12u
m7057 3687 3688 VSS VSS nch l=0.04u w=0.8u
m7058 3690 3689 VSS VSS nch l=0.04u w=0.8u
m7059 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m7060 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m7061 VSS 3722 3664 VSS nch l=0.04u w=0.4u
m7062 VSS 3452 VSS VSS nch l=0.26u w=0.8u
m7063 3680 3526 71434 VSS nch l=0.04u w=0.8u
m7064 VSS 3719 71435 VSS nch l=0.04u w=0.12u
m7065 3673 4351 71436 VSS nch l=0.04u w=0.8u
m7066 71441 3644 VSS VSS nch l=0.04u w=0.8u
m7067 71442 3645 VSS VSS nch l=0.04u w=0.8u
m7068 71443 3646 VSS VSS nch l=0.04u w=0.8u
m7069 71444 3647 VSS VSS nch l=0.04u w=0.8u
m7070 71445 3648 VSS VSS nch l=0.04u w=0.8u
m7071 71446 3649 VSS VSS nch l=0.04u w=0.8u
m7072 71447 3650 VSS VSS nch l=0.04u w=0.8u
m7073 71448 3651 VSS VSS nch l=0.04u w=0.8u
m7074 71449 3652 VSS VSS nch l=0.04u w=0.8u
m7075 71450 3653 VSS VSS nch l=0.04u w=0.8u
m7076 71451 3764 VSS VSS nch l=0.04u w=0.8u
m7077 3708 4062 VSS VSS nch l=0.04u w=0.4u
m7078 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m7079 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m7080 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m7081 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m7082 VSS 3612 71437 VSS nch l=0.04u w=0.12u
m7083 VSS 3611 71438 VSS nch l=0.04u w=0.12u
m7084 VSS 3614 71439 VSS nch l=0.04u w=0.12u
m7085 VSS 3613 71440 VSS nch l=0.04u w=0.12u
m7086 71452 3664 VSS VSS nch l=0.04u w=0.12u
m7087 3712 3711 VSS VSS nch l=0.04u w=0.8u
m7088 VSS 3692 3692 VSS nch l=0.04u w=0.8u
m7089 71453 3636 VSS VSS nch l=0.04u w=0.8u
m7090 71454 2508 VSS VSS nch l=0.04u w=0.8u
m7091 3719 3667 VSS VSS nch l=0.04u w=0.4u
m7092 3715 4328 3681 VSS nch l=0.04u w=0.4u
m7093 3716 4328 3682 VSS nch l=0.04u w=0.4u
m7094 71455 3478 3693 VSS nch l=0.04u w=0.8u
m7095 3694 3539 71441 VSS nch l=0.04u w=0.8u
m7096 71456 3483 3695 VSS nch l=0.04u w=0.8u
m7097 3696 3540 71442 VSS nch l=0.04u w=0.8u
m7098 3717 4328 3683 VSS nch l=0.04u w=0.4u
m7099 3718 4328 3684 VSS nch l=0.04u w=0.4u
m7100 71457 3479 3697 VSS nch l=0.04u w=0.8u
m7101 3698 3543 71443 VSS nch l=0.04u w=0.8u
m7102 3699 3544 71444 VSS nch l=0.04u w=0.8u
m7103 3700 3545 71445 VSS nch l=0.04u w=0.8u
m7104 71458 3201 3701 VSS nch l=0.04u w=0.8u
m7105 3702 3546 71446 VSS nch l=0.04u w=0.8u
m7106 3703 3547 71447 VSS nch l=0.04u w=0.8u
m7107 3704 3548 71448 VSS nch l=0.04u w=0.8u
m7108 71459 3202 3705 VSS nch l=0.04u w=0.8u
m7109 3706 3549 71449 VSS nch l=0.04u w=0.8u
m7110 3707 3550 71450 VSS nch l=0.04u w=0.8u
m7111 3642 3800 71451 VSS nch l=0.04u w=0.8u
m7112 3720 3685 3662 VSS nch l=0.04u w=0.4u
m7113 3721 3686 3663 VSS nch l=0.04u w=0.4u
m7114 3612 3674 VSS VSS nch l=0.04u w=0.4u
m7115 3611 3675 VSS VSS nch l=0.04u w=0.4u
m7116 3614 3676 VSS VSS nch l=0.04u w=0.4u
m7117 3613 3677 VSS VSS nch l=0.04u w=0.4u
m7118 VSS 3487 VSS VSS nch l=0.26u w=0.8u
m7119 VSS 3488 VSS VSS nch l=0.26u w=0.8u
m7120 3722 4251 71452 VSS nch l=0.04u w=0.12u
m7121 VSS 3709 3709 VSS nch l=0.04u w=0.8u
m7122 3713 3566 71453 VSS nch l=0.04u w=0.8u
m7123 3714 3180 71454 VSS nch l=0.04u w=0.8u
m7124 3725 3569 VSS VSS nch l=0.04u w=0.4u
m7125 71461 3624 3715 VSS nch l=0.04u w=0.12u
m7126 71462 3625 3716 VSS nch l=0.04u w=0.12u
m7127 VSS 3479 71455 VSS nch l=0.04u w=0.8u
m7128 VSS 1998 71456 VSS nch l=0.04u w=0.8u
m7129 71463 3626 3717 VSS nch l=0.04u w=0.12u
m7130 71464 3627 3718 VSS nch l=0.04u w=0.12u
m7131 VSS FRAC[13] 71457 VSS nch l=0.04u w=0.8u
m7132 VSS 3087 71458 VSS nch l=0.04u w=0.8u
m7133 VSS FRAC[13] 71459 VSS nch l=0.04u w=0.8u
m7134 71465 3800 3642 VSS nch l=0.04u w=0.8u
m7135 3726 3673 VSS VSS nch l=0.04u w=0.4u
m7136 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m7137 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m7138 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m7139 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m7140 71466 4062 VSS VSS nch l=0.04u w=0.8u
m7141 71467 4328 3720 VSS nch l=0.04u w=0.12u
m7142 71468 4328 3721 VSS nch l=0.04u w=0.12u
m7143 3728 3729 VSS VSS nch l=0.04u w=0.8u
m7144 3731 3730 VSS VSS nch l=0.04u w=0.8u
m7145 3732 3756 3722 VSS nch l=0.04u w=0.4u
m7146 VSS 3691 VSS VSS nch l=0.26u w=0.8u
m7147 VSS 3724 3724 VSS nch l=0.04u w=0.8u
m7148 71471 2445 VSS VSS nch l=0.04u w=0.8u
m7149 3736 3401 3725 VSS nch l=0.04u w=0.4u
m7150 VSS 3759 71461 VSS nch l=0.04u w=0.12u
m7151 VSS 3608 71462 VSS nch l=0.04u w=0.12u
m7152 VSS 3760 71463 VSS nch l=0.04u w=0.12u
m7153 VSS 3610 71464 VSS nch l=0.04u w=0.12u
m7154 VSS 3764 71465 VSS nch l=0.04u w=0.8u
m7155 3738 3592 VSS VSS nch l=0.04u w=0.4u
m7156 3740 3594 VSS VSS nch l=0.04u w=0.4u
m7157 3742 3596 VSS VSS nch l=0.04u w=0.4u
m7158 3743 3598 VSS VSS nch l=0.04u w=0.4u
m7159 3744 3599 VSS VSS nch l=0.04u w=0.4u
m7160 3746 3601 VSS VSS nch l=0.04u w=0.4u
m7161 3747 3602 VSS VSS nch l=0.04u w=0.4u
m7162 3748 3603 VSS VSS nch l=0.04u w=0.4u
m7163 3750 3605 VSS VSS nch l=0.04u w=0.4u
m7164 3751 3606 VSS VSS nch l=0.04u w=0.4u
m7165 3727 2245 71466 VSS nch l=0.04u w=0.8u
m7166 VSS 3766 71467 VSS nch l=0.04u w=0.12u
m7167 VSS 3767 71468 VSS nch l=0.04u w=0.12u
m7168 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7169 VSS 3733 3733 VSS nch l=0.04u w=0.8u
m7170 71477 3713 VSS VSS nch l=0.04u w=0.8u
m7171 3735 3180 71471 VSS nch l=0.04u w=0.8u
m7172 3758 3180 VSS VSS nch l=0.04u w=0.4u
m7173 3401 3725 3736 VSS nch l=0.04u w=0.4u
m7174 3759 3715 VSS VSS nch l=0.04u w=0.4u
m7175 3608 3716 VSS VSS nch l=0.04u w=0.4u
m7176 VSS 3529 VSS VSS nch l=0.26u w=0.8u
m7177 VSS 3530 VSS VSS nch l=0.26u w=0.8u
m7178 3760 3717 VSS VSS nch l=0.04u w=0.4u
m7179 3610 3718 VSS VSS nch l=0.04u w=0.4u
m7180 VSS 3533 VSS VSS nch l=0.26u w=0.8u
m7181 VSS 3534 VSS VSS nch l=0.26u w=0.8u
m7182 3633 3413 3738 VSS nch l=0.04u w=0.4u
m7183 3762 3415 3740 VSS nch l=0.04u w=0.4u
m7184 3609 3417 3742 VSS nch l=0.04u w=0.4u
m7185 3582 3418 3743 VSS nch l=0.04u w=0.4u
m7186 3587 3419 3744 VSS nch l=0.04u w=0.4u
m7187 3586 3421 3746 VSS nch l=0.04u w=0.4u
m7188 3622 3422 3747 VSS nch l=0.04u w=0.4u
m7189 3589 3423 3748 VSS nch l=0.04u w=0.4u
m7190 3588 3425 3750 VSS nch l=0.04u w=0.4u
m7191 3623 3426 3751 VSS nch l=0.04u w=0.4u
m7192 71482 3726 VSS VSS nch l=0.04u w=0.8u
m7193 3766 3720 VSS VSS nch l=0.04u w=0.4u
m7194 3767 3721 VSS VSS nch l=0.04u w=0.4u
m7195 VSS 3752 3752 VSS nch l=0.04u w=0.8u
m7196 VSS 3755 3755 VSS nch l=0.04u w=0.8u
m7197 VSS 3691 VSS VSS nch l=0.26u w=0.8u
m7198 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7199 VSS 4251 3756 VSS nch l=0.04u w=0.4u
m7200 3757 3665 71477 VSS nch l=0.04u w=0.8u
m7201 3768 2508 3758 VSS nch l=0.04u w=0.4u
m7202 3769 3770 VSS VSS nch l=0.04u w=0.8u
m7203 3772 3771 VSS VSS nch l=0.04u w=0.8u
m7204 3773 3774 VSS VSS nch l=0.04u w=0.8u
m7205 3776 3775 VSS VSS nch l=0.04u w=0.8u
m7206 3413 3738 3633 VSS nch l=0.04u w=0.4u
m7207 3415 3740 3762 VSS nch l=0.04u w=0.4u
m7208 3417 3742 3609 VSS nch l=0.04u w=0.4u
m7209 3418 3743 3582 VSS nch l=0.04u w=0.4u
m7210 3419 3744 3587 VSS nch l=0.04u w=0.4u
m7211 3421 3746 3586 VSS nch l=0.04u w=0.4u
m7212 3422 3747 3622 VSS nch l=0.04u w=0.4u
m7213 3423 3748 3589 VSS nch l=0.04u w=0.4u
m7214 3425 3750 3588 VSS nch l=0.04u w=0.4u
m7215 3426 3751 3623 VSS nch l=0.04u w=0.4u
m7216 71483 3862 3764 VSS nch l=0.04u w=0.8u
m7217 71484 3643 71482 VSS nch l=0.04u w=0.8u
m7218 3632 3784 3737 VSS nch l=0.04u w=0.4u
m7219 3761 3785 3739 VSS nch l=0.04u w=0.4u
m7220 3763 3786 3741 VSS nch l=0.04u w=0.4u
m7221 3407 3791 3745 VSS nch l=0.04u w=0.4u
m7222 3409 3796 3749 VSS nch l=0.04u w=0.4u
m7223 71490 3708 VSS VSS nch l=0.04u w=0.8u
m7224 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7225 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7226 71491 3665 3757 VSS nch l=0.04u w=0.8u
m7227 2508 3758 3768 VSS nch l=0.04u w=0.4u
m7228 3783 3735 VSS VSS nch l=0.04u w=0.4u
m7229 VSS 3835 71483 VSS nch l=0.04u w=0.8u
m7230 3765 3953 71484 VSS nch l=0.04u w=0.8u
m7231 3784 3737 3632 VSS nch l=0.04u w=0.4u
m7232 3785 3739 3761 VSS nch l=0.04u w=0.4u
m7233 3786 3741 3763 VSS nch l=0.04u w=0.4u
m7234 3791 3745 3407 VSS nch l=0.04u w=0.4u
m7235 3796 3749 3409 VSS nch l=0.04u w=0.4u
m7236 3782 3654 71490 VSS nch l=0.04u w=0.8u
m7237 3797 4328 3766 VSS nch l=0.04u w=0.4u
m7238 3798 4328 3767 VSS nch l=0.04u w=0.4u
m7239 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7240 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7241 VSS 3691 VSS VSS nch l=0.26u w=0.8u
m7242 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7243 71510 3846 VSS VSS nch l=0.04u w=0.8u
m7244 VSS 3713 71491 VSS nch l=0.04u w=0.8u
m7245 3799 3680 VSS VSS nch l=0.04u w=0.4u
m7246 VSS 3777 3784 VSS nch l=0.04u w=0.4u
m7247 VSS 3778 3785 VSS nch l=0.04u w=0.4u
m7248 VSS 3779 3786 VSS nch l=0.04u w=0.4u
m7249 VSS 3788 3788 VSS nch l=0.04u w=0.8u
m7250 VSS 3789 3789 VSS nch l=0.04u w=0.8u
m7251 VSS 3780 3791 VSS nch l=0.04u w=0.4u
m7252 VSS 3793 3793 VSS nch l=0.04u w=0.8u
m7253 VSS 3794 3794 VSS nch l=0.04u w=0.8u
m7254 VSS 3781 3796 VSS nch l=0.04u w=0.4u
m7255 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7256 71512 3685 3797 VSS nch l=0.04u w=0.12u
m7257 71513 3686 3798 VSS nch l=0.04u w=0.12u
m7258 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7259 3732 3867 71510 VSS nch l=0.04u w=0.8u
m7260 71514 1200 3800 VSS nch l=0.04u w=0.8u
m7261 3818 PD VSS VSS nch l=0.04u w=0.4u
m7262 3819 3694 VSS VSS nch l=0.04u w=0.4u
m7263 3820 3696 VSS VSS nch l=0.04u w=0.4u
m7264 3821 3698 VSS VSS nch l=0.04u w=0.4u
m7265 3822 3699 VSS VSS nch l=0.04u w=0.4u
m7266 3823 3700 VSS VSS nch l=0.04u w=0.4u
m7267 3824 3702 VSS VSS nch l=0.04u w=0.4u
m7268 3825 3703 VSS VSS nch l=0.04u w=0.4u
m7269 3826 3704 VSS VSS nch l=0.04u w=0.4u
m7270 3827 3706 VSS VSS nch l=0.04u w=0.4u
m7271 3828 3707 VSS VSS nch l=0.04u w=0.4u
m7272 71515 3782 VSS VSS nch l=0.04u w=0.8u
m7273 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7274 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7275 VSS 3833 71512 VSS nch l=0.04u w=0.12u
m7276 VSS 3834 71513 VSS nch l=0.04u w=0.12u
m7277 VSS 3691 VSS VSS nch l=0.26u w=0.8u
m7278 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7279 VSS 3801 3801 VSS nch l=0.04u w=0.8u
m7280 VSS 3804 3804 VSS nch l=0.04u w=0.8u
m7281 VSS 3805 3805 VSS nch l=0.04u w=0.8u
m7282 VSS 3808 3808 VSS nch l=0.04u w=0.8u
m7283 VSS 3809 3809 VSS nch l=0.04u w=0.8u
m7284 VSS 3812 3812 VSS nch l=0.04u w=0.8u
m7285 VSS 3813 3813 VSS nch l=0.04u w=0.8u
m7286 VSS 3816 3816 VSS nch l=0.04u w=0.8u
m7287 71516 3867 3732 VSS nch l=0.04u w=0.8u
m7288 3830 4251 VSS VSS nch l=0.04u w=0.4u
m7289 VSS 3787 VSS VSS nch l=0.26u w=0.8u
m7290 VSS 3790 VSS VSS nch l=0.26u w=0.8u
m7291 VSS 3792 VSS VSS nch l=0.26u w=0.8u
m7292 VSS 3795 VSS VSS nch l=0.26u w=0.8u
m7293 71517 3768 3817 VSS nch l=0.04u w=0.8u
m7294 VSS 4062 71514 VSS nch l=0.04u w=0.8u
m7295 71518 2761 VSS VSS nch l=0.04u w=0.8u
m7296 71519 3939 3455 VSS nch l=0.04u w=0.8u
m7297 71520 3940 3457 VSS nch l=0.04u w=0.8u
m7298 71521 3941 3459 VSS nch l=0.04u w=0.8u
m7299 71522 3942 3463 VSS nch l=0.04u w=0.8u
m7300 71523 3943 3467 VSS nch l=0.04u w=0.8u
m7301 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7302 3829 3727 71515 VSS nch l=0.04u w=0.8u
m7303 3833 3797 VSS VSS nch l=0.04u w=0.4u
m7304 3834 3798 VSS VSS nch l=0.04u w=0.4u
m7305 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7306 VSS 3846 71516 VSS nch l=0.04u w=0.8u
m7307 VSS 3666 71517 VSS nch l=0.04u w=0.8u
m7308 71525 3025 71518 VSS nch l=0.04u w=0.8u
m7309 VSS 3854 71519 VSS nch l=0.04u w=0.8u
m7310 VSS 3855 71520 VSS nch l=0.04u w=0.8u
m7311 VSS 3856 71521 VSS nch l=0.04u w=0.8u
m7312 VSS 3857 71522 VSS nch l=0.04u w=0.8u
m7313 VSS 3858 71523 VSS nch l=0.04u w=0.8u
m7314 VSS 4251 3832 VSS nch l=0.04u w=0.4u
m7315 71527 2780 VSS VSS nch l=0.04u w=0.8u
m7316 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7317 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7318 71528 2781 VSS VSS nch l=0.04u w=0.8u
m7319 71529 2782 VSS VSS nch l=0.04u w=0.8u
m7320 71530 2786 VSS VSS nch l=0.04u w=0.8u
m7321 71531 2787 VSS VSS nch l=0.04u w=0.8u
m7322 71532 2788 VSS VSS nch l=0.04u w=0.8u
m7323 71533 2789 VSS VSS nch l=0.04u w=0.8u
m7324 71534 2790 VSS VSS nch l=0.04u w=0.8u
m7325 71535 2791 VSS VSS nch l=0.04u w=0.8u
m7326 71536 2792 VSS VSS nch l=0.04u w=0.8u
m7327 71537 3727 3829 VSS nch l=0.04u w=0.8u
m7328 VSS 3691 VSS VSS nch l=0.26u w=0.8u
m7329 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7330 VSS 3802 VSS VSS nch l=0.26u w=0.8u
m7331 VSS 3803 VSS VSS nch l=0.26u w=0.8u
m7332 VSS 3806 VSS VSS nch l=0.26u w=0.8u
m7333 VSS 3807 VSS VSS nch l=0.26u w=0.8u
m7334 VSS 3810 VSS VSS nch l=0.26u w=0.8u
m7335 VSS 3811 VSS VSS nch l=0.26u w=0.8u
m7336 VSS 3814 VSS VSS nch l=0.26u w=0.8u
m7337 VSS 3815 VSS VSS nch l=0.26u w=0.8u
m7338 VSS 3787 VSS VSS nch l=0.26u w=0.8u
m7339 VSS 3790 VSS VSS nch l=0.26u w=0.8u
m7340 VSS 3792 VSS VSS nch l=0.26u w=0.8u
m7341 VSS 3795 VSS VSS nch l=0.26u w=0.8u
m7342 3847 3830 3757 VSS nch l=0.04u w=0.4u
m7343 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7344 3831 3302 71525 VSS nch l=0.04u w=0.8u
m7345 VSS 4062 3835 VSS nch l=0.04u w=0.4u
m7346 71538 3047 71527 VSS nch l=0.04u w=0.8u
m7347 71539 3049 71528 VSS nch l=0.04u w=0.8u
m7348 71540 3051 71529 VSS nch l=0.04u w=0.8u
m7349 71541 3053 71530 VSS nch l=0.04u w=0.8u
m7350 71542 3054 71531 VSS nch l=0.04u w=0.8u
m7351 71543 3056 71532 VSS nch l=0.04u w=0.8u
m7352 71544 3057 71533 VSS nch l=0.04u w=0.8u
m7353 71545 3058 71534 VSS nch l=0.04u w=0.8u
m7354 71546 3060 71535 VSS nch l=0.04u w=0.8u
m7355 71547 3061 71536 VSS nch l=0.04u w=0.8u
m7356 VSS 3782 71537 VSS nch l=0.04u w=0.8u
m7357 3849 3848 VSS VSS nch l=0.04u w=0.8u
m7358 3850 4328 VSS VSS nch l=0.04u w=0.4u
m7359 3851 4328 VSS VSS nch l=0.04u w=0.4u
m7360 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7361 71548 3944 3846 VSS nch l=0.04u w=0.8u
m7362 71549 4251 3847 VSS nch l=0.04u w=0.12u
m7363 71550 3817 VSS VSS nch l=0.04u w=0.8u
m7364 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7365 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7366 71552 3737 VSS VSS nch l=0.04u w=0.8u
m7367 3836 3321 71538 VSS nch l=0.04u w=0.8u
m7368 71553 3739 VSS VSS nch l=0.04u w=0.8u
m7369 3837 3323 71539 VSS nch l=0.04u w=0.8u
m7370 71554 3741 VSS VSS nch l=0.04u w=0.8u
m7371 3838 3325 71540 VSS nch l=0.04u w=0.8u
m7372 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7373 3839 3327 71541 VSS nch l=0.04u w=0.8u
m7374 3840 3328 71542 VSS nch l=0.04u w=0.8u
m7375 71555 3745 VSS VSS nch l=0.04u w=0.8u
m7376 3841 3330 71543 VSS nch l=0.04u w=0.8u
m7377 3842 3331 71544 VSS nch l=0.04u w=0.8u
m7378 3843 3332 71545 VSS nch l=0.04u w=0.8u
m7379 71556 3749 VSS VSS nch l=0.04u w=0.8u
m7380 3844 3334 71546 VSS nch l=0.04u w=0.8u
m7381 3845 3335 71547 VSS nch l=0.04u w=0.8u
m7382 3853 3832 3765 VSS nch l=0.04u w=0.4u
m7383 VSS 3802 VSS VSS nch l=0.26u w=0.8u
m7384 VSS 3803 VSS VSS nch l=0.26u w=0.8u
m7385 VSS 3806 VSS VSS nch l=0.26u w=0.8u
m7386 VSS 3807 VSS VSS nch l=0.26u w=0.8u
m7387 VSS 3810 VSS VSS nch l=0.26u w=0.8u
m7388 VSS 3811 VSS VSS nch l=0.26u w=0.8u
m7389 VSS 3814 VSS VSS nch l=0.26u w=0.8u
m7390 VSS 3815 VSS VSS nch l=0.26u w=0.8u
m7391 VSS 3899 71548 VSS nch l=0.04u w=0.8u
m7392 VSS 3787 VSS VSS nch l=0.26u w=0.8u
m7393 VSS 3790 VSS VSS nch l=0.26u w=0.8u
m7394 VSS 3792 VSS VSS nch l=0.26u w=0.8u
m7395 VSS 3795 VSS VSS nch l=0.26u w=0.8u
m7396 VSS 3868 71549 VSS nch l=0.04u w=0.12u
m7397 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7398 3852 3714 71550 VSS nch l=0.04u w=0.8u
m7399 3861 3831 VSS VSS nch l=0.04u w=0.4u
m7400 3854 3777 71552 VSS nch l=0.04u w=0.8u
m7401 3855 3778 71553 VSS nch l=0.04u w=0.8u
m7402 3856 3779 71554 VSS nch l=0.04u w=0.8u
m7403 3857 3780 71555 VSS nch l=0.04u w=0.8u
m7404 3858 3781 71556 VSS nch l=0.04u w=0.8u
m7405 3862 3869 3518 VSS nch l=0.04u w=0.4u
m7406 71558 4251 3853 VSS nch l=0.04u w=0.24u
m7407 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7408 3863 4251 VSS VSS nch l=0.04u w=0.4u
m7409 VSS 3860 3860 VSS nch l=0.04u w=0.8u
m7410 3864 3850 3833 VSS nch l=0.04u w=0.4u
m7411 3865 3851 3834 VSS nch l=0.04u w=0.4u
m7412 3868 3847 VSS VSS nch l=0.04u w=0.4u
m7413 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7414 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7415 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7416 VSS 3802 VSS VSS nch l=0.26u w=0.8u
m7417 VSS 3803 VSS VSS nch l=0.26u w=0.8u
m7418 VSS 3806 VSS VSS nch l=0.26u w=0.8u
m7419 VSS 3807 VSS VSS nch l=0.26u w=0.8u
m7420 VSS 3810 VSS VSS nch l=0.26u w=0.8u
m7421 VSS 3811 VSS VSS nch l=0.26u w=0.8u
m7422 VSS 3814 VSS VSS nch l=0.26u w=0.8u
m7423 VSS 3815 VSS VSS nch l=0.26u w=0.8u
m7424 3869 3518 3862 VSS nch l=0.04u w=0.4u
m7425 VSS 3881 71558 VSS nch l=0.04u w=0.24u
m7426 3870 3836 VSS VSS nch l=0.04u w=0.4u
m7427 3871 3837 VSS VSS nch l=0.04u w=0.4u
m7428 3872 3838 VSS VSS nch l=0.04u w=0.4u
m7429 3873 3839 VSS VSS nch l=0.04u w=0.4u
m7430 3874 3840 VSS VSS nch l=0.04u w=0.4u
m7431 3875 3841 VSS VSS nch l=0.04u w=0.4u
m7432 3876 3842 VSS VSS nch l=0.04u w=0.4u
m7433 3877 3843 VSS VSS nch l=0.04u w=0.4u
m7434 3878 3844 VSS VSS nch l=0.04u w=0.4u
m7435 3879 3845 VSS VSS nch l=0.04u w=0.4u
m7436 71560 4328 3864 VSS nch l=0.04u w=0.12u
m7437 71561 4328 3865 VSS nch l=0.04u w=0.12u
m7438 VSS 3787 VSS VSS nch l=0.26u w=0.8u
m7439 VSS 3790 VSS VSS nch l=0.26u w=0.8u
m7440 VSS 3792 VSS VSS nch l=0.26u w=0.8u
m7441 VSS 3795 VSS VSS nch l=0.26u w=0.8u
m7442 71567 FBDIV[9] 3867 VSS nch l=0.04u w=0.8u
m7443 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7444 3880 3768 VSS VSS nch l=0.04u w=0.4u
m7445 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7446 71568 3818 VSS VSS nch l=0.04u w=0.8u
m7447 VSS 3859 VSS VSS nch l=0.26u w=0.8u
m7448 71569 3861 VSS VSS nch l=0.04u w=0.8u
m7449 3884 3863 3829 VSS nch l=0.04u w=0.4u
m7450 VSS 3897 71560 VSS nch l=0.04u w=0.12u
m7451 VSS 3898 71561 VSS nch l=0.04u w=0.12u
m7452 VSS 4062 71567 VSS nch l=0.04u w=0.8u
m7453 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7454 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7455 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7456 3885 4251 3868 VSS nch l=0.04u w=0.4u
m7457 VSS 3802 VSS VSS nch l=0.26u w=0.8u
m7458 VSS 3803 VSS VSS nch l=0.26u w=0.8u
m7459 VSS 3806 VSS VSS nch l=0.26u w=0.8u
m7460 VSS 3807 VSS VSS nch l=0.26u w=0.8u
m7461 VSS 3810 VSS VSS nch l=0.26u w=0.8u
m7462 VSS 3811 VSS VSS nch l=0.26u w=0.8u
m7463 VSS 3814 VSS VSS nch l=0.26u w=0.8u
m7464 VSS 3815 VSS VSS nch l=0.26u w=0.8u
m7465 3886 3666 3880 VSS nch l=0.04u w=0.4u
m7466 3881 3853 71568 VSS nch l=0.04u w=0.8u
m7467 71573 3569 71569 VSS nch l=0.04u w=0.8u
m7468 VSS 3869 3883 VSS nch l=0.04u w=0.4u
m7469 3777 3900 3760 VSS nch l=0.04u w=0.4u
m7470 71574 3870 VSS VSS nch l=0.04u w=0.8u
m7471 3778 3901 1963 VSS nch l=0.04u w=0.4u
m7472 71575 3871 VSS VSS nch l=0.04u w=0.8u
m7473 3779 3902 FRAC[12] VSS nch l=0.04u w=0.4u
m7474 71576 3872 VSS VSS nch l=0.04u w=0.8u
m7475 71577 3873 VSS VSS nch l=0.04u w=0.8u
m7476 71578 3874 VSS VSS nch l=0.04u w=0.8u
m7477 3780 3903 3409 VSS nch l=0.04u w=0.4u
m7478 71579 3875 VSS VSS nch l=0.04u w=0.8u
m7479 71580 3876 VSS VSS nch l=0.04u w=0.8u
m7480 71581 3877 VSS VSS nch l=0.04u w=0.8u
m7481 3781 3904 FRAC[12] VSS nch l=0.04u w=0.4u
m7482 71582 3878 VSS VSS nch l=0.04u w=0.8u
m7483 71583 3879 VSS VSS nch l=0.04u w=0.8u
m7484 71584 4251 3884 VSS nch l=0.04u w=0.12u
m7485 3897 3864 VSS VSS nch l=0.04u w=0.4u
m7486 3898 3865 VSS VSS nch l=0.04u w=0.4u
m7487 VSS 3787 VSS VSS nch l=0.26u w=0.8u
m7488 VSS 3790 VSS VSS nch l=0.26u w=0.8u
m7489 VSS 3792 VSS VSS nch l=0.26u w=0.8u
m7490 VSS 3795 VSS VSS nch l=0.26u w=0.8u
m7491 VSS 3710 VSS VSS nch l=0.26u w=0.8u
m7492 71587 3830 3885 VSS nch l=0.04u w=0.12u
m7493 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7494 VSS 3859 VSS VSS nch l=0.26u w=0.8u
m7495 3666 3880 3886 VSS nch l=0.04u w=0.4u
m7496 3882 2667 71573 VSS nch l=0.04u w=0.8u
m7497 3900 3760 3777 VSS nch l=0.04u w=0.4u
m7498 71588 3592 71574 VSS nch l=0.04u w=0.8u
m7499 3901 1963 3778 VSS nch l=0.04u w=0.4u
m7500 71589 3594 71575 VSS nch l=0.04u w=0.8u
m7501 3902 FRAC[12] 3779 VSS nch l=0.04u w=0.4u
m7502 71590 3596 71576 VSS nch l=0.04u w=0.8u
m7503 71591 3598 71577 VSS nch l=0.04u w=0.8u
m7504 71592 3599 71578 VSS nch l=0.04u w=0.8u
m7505 3903 3409 3780 VSS nch l=0.04u w=0.4u
m7506 71593 3601 71579 VSS nch l=0.04u w=0.8u
m7507 71594 3602 71580 VSS nch l=0.04u w=0.8u
m7508 71595 3603 71581 VSS nch l=0.04u w=0.8u
m7509 3904 FRAC[12] 3781 VSS nch l=0.04u w=0.4u
m7510 71596 3605 71582 VSS nch l=0.04u w=0.8u
m7511 71597 3606 71583 VSS nch l=0.04u w=0.8u
m7512 VSS 3916 71584 VSS nch l=0.04u w=0.12u
m7513 3906 3905 VSS VSS nch l=0.04u w=0.8u
m7514 3907 3908 VSS VSS nch l=0.04u w=0.8u
m7515 3910 3909 VSS VSS nch l=0.04u w=0.8u
m7516 3911 3912 VSS VSS nch l=0.04u w=0.8u
m7517 3913 3914 VSS VSS nch l=0.04u w=0.8u
m7518 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7519 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7520 VSS 4062 3899 VSS nch l=0.04u w=0.4u
m7521 VSS 3723 VSS VSS nch l=0.26u w=0.8u
m7522 VSS 3802 VSS VSS nch l=0.26u w=0.8u
m7523 VSS 3803 VSS VSS nch l=0.26u w=0.8u
m7524 VSS 3806 VSS VSS nch l=0.26u w=0.8u
m7525 VSS 3807 VSS VSS nch l=0.26u w=0.8u
m7526 VSS 3810 VSS VSS nch l=0.26u w=0.8u
m7527 VSS 3811 VSS VSS nch l=0.26u w=0.8u
m7528 VSS 3814 VSS VSS nch l=0.26u w=0.8u
m7529 VSS 3815 VSS VSS nch l=0.26u w=0.8u
m7530 VSS 3590 71587 VSS nch l=0.04u w=0.12u
m7531 3915 4251 3881 VSS nch l=0.04u w=0.4u
m7532 VSS 3759 3900 VSS nch l=0.04u w=0.4u
m7533 3887 2678 71588 VSS nch l=0.04u w=0.8u
m7534 VSS 3763 3901 VSS nch l=0.04u w=0.4u
m7535 3888 2679 71589 VSS nch l=0.04u w=0.8u
m7536 VSS 3760 3902 VSS nch l=0.04u w=0.4u
m7537 3889 2680 71590 VSS nch l=0.04u w=0.8u
m7538 3890 2683 71591 VSS nch l=0.04u w=0.8u
m7539 3891 2684 71592 VSS nch l=0.04u w=0.8u
m7540 VSS 3553 3903 VSS nch l=0.04u w=0.4u
m7541 3892 2685 71593 VSS nch l=0.04u w=0.8u
m7542 3893 2686 71594 VSS nch l=0.04u w=0.8u
m7543 3894 2687 71595 VSS nch l=0.04u w=0.8u
m7544 VSS 3554 3904 VSS nch l=0.04u w=0.4u
m7545 3895 2688 71596 VSS nch l=0.04u w=0.8u
m7546 3896 2689 71597 VSS nch l=0.04u w=0.8u
m7547 VSS 3953 3869 VSS nch l=0.04u w=0.4u
m7548 3916 3884 VSS VSS nch l=0.04u w=0.4u
m7549 3917 4328 3897 VSS nch l=0.04u w=0.4u
m7550 3918 4328 3898 VSS nch l=0.04u w=0.4u
m7551 3920 3919 VSS VSS nch l=0.04u w=0.8u
m7552 3921 3922 VSS VSS nch l=0.04u w=0.8u
m7553 3924 3923 VSS VSS nch l=0.04u w=0.8u
m7554 3925 3926 VSS VSS nch l=0.04u w=0.8u
m7555 3928 3927 VSS VSS nch l=0.04u w=0.8u
m7556 3929 3930 VSS VSS nch l=0.04u w=0.8u
m7557 3932 3931 VSS VSS nch l=0.04u w=0.8u
m7558 3933 3934 VSS VSS nch l=0.04u w=0.8u
m7559 3936 3935 VSS VSS nch l=0.04u w=0.8u
m7560 VSS 3734 VSS VSS nch l=0.26u w=0.8u
m7561 3590 3885 VSS VSS nch l=0.04u w=0.4u
m7562 VSS 3859 VSS VSS nch l=0.26u w=0.8u
m7563 71604 3832 3915 VSS nch l=0.04u w=0.12u
m7564 3937 2445 VSS VSS nch l=0.04u w=0.4u
m7565 71605 3799 VSS VSS nch l=0.04u w=0.8u
m7566 71606 3850 3917 VSS nch l=0.04u w=0.12u
m7567 71607 3851 3918 VSS nch l=0.04u w=0.12u
m7568 VSS 3753 VSS VSS nch l=0.26u w=0.8u
m7569 VSS 3754 VSS VSS nch l=0.26u w=0.8u
m7570 3944 3958 3619 VSS nch l=0.04u w=0.4u
m7571 3945 3946 VSS VSS nch l=0.04u w=0.8u
m7572 VSS 4044 71604 VSS nch l=0.04u w=0.12u
m7573 VSS 3886 3937 VSS nch l=0.04u w=0.4u
m7574 3938 3882 71605 VSS nch l=0.04u w=0.8u
m7575 71611 3759 3939 VSS nch l=0.04u w=0.8u
m7576 71612 3819 VSS VSS nch l=0.04u w=0.8u
m7577 71613 3763 3940 VSS nch l=0.04u w=0.8u
m7578 71614 3820 VSS VSS nch l=0.04u w=0.8u
m7579 71615 3760 3941 VSS nch l=0.04u w=0.8u
m7580 71616 3821 VSS VSS nch l=0.04u w=0.8u
m7581 71617 3822 VSS VSS nch l=0.04u w=0.8u
m7582 71618 3823 VSS VSS nch l=0.04u w=0.8u
m7583 71619 3553 3942 VSS nch l=0.04u w=0.8u
m7584 71620 3824 VSS VSS nch l=0.04u w=0.8u
m7585 71621 3825 VSS VSS nch l=0.04u w=0.8u
m7586 71622 3826 VSS VSS nch l=0.04u w=0.8u
m7587 71623 3554 3943 VSS nch l=0.04u w=0.8u
m7588 71624 3827 VSS VSS nch l=0.04u w=0.8u
m7589 71625 3828 VSS VSS nch l=0.04u w=0.8u
m7590 3953 3963 VSS VSS nch l=0.04u w=0.4u
m7591 3947 4251 3916 VSS nch l=0.04u w=0.4u
m7592 VSS 2131 71606 VSS nch l=0.04u w=0.12u
m7593 VSS 3961 71607 VSS nch l=0.04u w=0.12u
m7594 3954 3955 VSS VSS nch l=0.04u w=0.8u
m7595 3957 3956 VSS VSS nch l=0.04u w=0.8u
m7596 3958 3619 3944 VSS nch l=0.04u w=0.4u
m7597 VSS 3859 VSS VSS nch l=0.26u w=0.8u
m7598 3959 3590 VSS VSS nch l=0.04u w=0.4u
m7599 3960 3915 VSS VSS nch l=0.04u w=0.4u
m7600 VSS 3760 71611 VSS nch l=0.04u w=0.8u
m7601 3737 3887 71612 VSS nch l=0.04u w=0.8u
m7602 VSS 1963 71613 VSS nch l=0.04u w=0.8u
m7603 3739 3888 71614 VSS nch l=0.04u w=0.8u
m7604 VSS FRAC[12] 71615 VSS nch l=0.04u w=0.8u
m7605 3741 3889 71616 VSS nch l=0.04u w=0.8u
m7606 3948 3890 71617 VSS nch l=0.04u w=0.8u
m7607 3949 3891 71618 VSS nch l=0.04u w=0.8u
m7608 VSS 3409 71619 VSS nch l=0.04u w=0.8u
m7609 3745 3892 71620 VSS nch l=0.04u w=0.8u
m7610 3950 3893 71621 VSS nch l=0.04u w=0.8u
m7611 3951 3894 71622 VSS nch l=0.04u w=0.8u
m7612 VSS FRAC[12] 71623 VSS nch l=0.04u w=0.8u
m7613 3749 3895 71624 VSS nch l=0.04u w=0.8u
m7614 3952 3896 71625 VSS nch l=0.04u w=0.8u
m7615 VSS 3963 3953 VSS nch l=0.04u w=0.4u
m7616 71629 3863 3947 VSS nch l=0.04u w=0.12u
m7617 2131 3917 VSS VSS nch l=0.04u w=0.4u
m7618 3961 3918 VSS VSS nch l=0.04u w=0.4u
m7619 VSS 3590 3959 VSS nch l=0.04u w=0.4u
m7620 VSS 3661 71629 VSS nch l=0.04u w=0.12u
m7621 VSS 3859 VSS VSS nch l=0.26u w=0.8u
m7622 VSS 3958 3962 VSS nch l=0.04u w=0.4u
m7623 71656 3818 VSS VSS nch l=0.04u w=0.8u
m7624 3661 3947 VSS VSS nch l=0.04u w=0.4u
m7625 VSS 4042 3963 VSS nch l=0.04u w=0.4u
m7626 3965 2131 VSS VSS nch l=0.04u w=0.4u
m7627 3966 4328 VSS VSS nch l=0.04u w=0.4u
m7628 3968 3967 VSS VSS nch l=0.04u w=0.8u
m7629 3969 3959 VSS VSS nch l=0.04u w=0.4u
m7630 3964 3960 71656 VSS nch l=0.04u w=0.8u
m7631 71693 3963 VSS VSS nch l=0.04u w=0.12u
m7632 71696 3953 3958 VSS nch l=0.04u w=0.8u
m7633 4042 4059 71693 VSS nch l=0.04u w=0.12u
m7634 4040 3661 VSS VSS nch l=0.04u w=0.4u
m7635 VSS 3970 3970 VSS nch l=0.04u w=0.8u
m7636 VSS 3973 3973 VSS nch l=0.04u w=0.8u
m7637 VSS 3974 3974 VSS nch l=0.04u w=0.8u
m7638 VSS 3977 3977 VSS nch l=0.04u w=0.8u
m7639 VSS 3978 3978 VSS nch l=0.04u w=0.8u
m7640 VSS 3981 3981 VSS nch l=0.04u w=0.8u
m7641 VSS 3982 3982 VSS nch l=0.04u w=0.8u
m7642 VSS 3985 3985 VSS nch l=0.04u w=0.8u
m7643 VSS 3986 3986 VSS nch l=0.04u w=0.8u
m7644 VSS 3989 3989 VSS nch l=0.04u w=0.8u
m7645 VSS 3990 3990 VSS nch l=0.04u w=0.8u
m7646 VSS 3993 3993 VSS nch l=0.04u w=0.8u
m7647 VSS 3994 3994 VSS nch l=0.04u w=0.8u
m7648 VSS 3997 3997 VSS nch l=0.04u w=0.8u
m7649 VSS 3998 3998 VSS nch l=0.04u w=0.8u
m7650 VSS 4001 4001 VSS nch l=0.04u w=0.8u
m7651 VSS 4002 4002 VSS nch l=0.04u w=0.8u
m7652 VSS 4005 4005 VSS nch l=0.04u w=0.8u
m7653 VSS 4006 4006 VSS nch l=0.04u w=0.8u
m7654 VSS 4009 4009 VSS nch l=0.04u w=0.8u
m7655 4043 4230 VSS VSS nch l=0.04u w=0.4u
m7656 4041 3966 3961 VSS nch l=0.04u w=0.4u
m7657 VSS 4010 4010 VSS nch l=0.04u w=0.8u
m7658 VSS 4013 4013 VSS nch l=0.04u w=0.8u
m7659 VSS 4014 4014 VSS nch l=0.04u w=0.8u
m7660 VSS 4017 4017 VSS nch l=0.04u w=0.8u
m7661 VSS 4018 4018 VSS nch l=0.04u w=0.8u
m7662 VSS 4021 4021 VSS nch l=0.04u w=0.8u
m7663 VSS 4022 4022 VSS nch l=0.04u w=0.8u
m7664 VSS 4025 4025 VSS nch l=0.04u w=0.8u
m7665 VSS 4026 4026 VSS nch l=0.04u w=0.8u
m7666 VSS 4029 4029 VSS nch l=0.04u w=0.8u
m7667 VSS 4030 4030 VSS nch l=0.04u w=0.8u
m7668 VSS 4033 4033 VSS nch l=0.04u w=0.8u
m7669 VSS 4034 4034 VSS nch l=0.04u w=0.8u
m7670 VSS 4037 4037 VSS nch l=0.04u w=0.8u
m7671 VSS 4039 4039 VSS nch l=0.04u w=0.8u
m7672 VSS 4048 71696 VSS nch l=0.04u w=0.8u
m7673 71699 3524 VSS VSS nch l=0.04u w=0.8u
m7674 4044 3964 VSS VSS nch l=0.04u w=0.4u
m7675 4045 4251 4042 VSS nch l=0.04u w=0.4u
m7676 VSS 3661 4040 VSS nch l=0.04u w=0.4u
m7677 71700 4328 4041 VSS nch l=0.04u w=0.12u
m7678 4047 4328 VSS VSS nch l=0.04u w=0.4u
m7679 3567 3969 71699 VSS nch l=0.04u w=0.8u
m7680 VSS 3971 VSS VSS nch l=0.26u w=0.8u
m7681 VSS 3972 VSS VSS nch l=0.26u w=0.8u
m7682 VSS 3975 VSS VSS nch l=0.26u w=0.8u
m7683 VSS 3976 VSS VSS nch l=0.26u w=0.8u
m7684 VSS 3979 VSS VSS nch l=0.26u w=0.8u
m7685 VSS 3980 VSS VSS nch l=0.26u w=0.8u
m7686 VSS 3983 VSS VSS nch l=0.26u w=0.8u
m7687 VSS 3984 VSS VSS nch l=0.26u w=0.8u
m7688 VSS 3987 VSS VSS nch l=0.26u w=0.8u
m7689 VSS 3988 VSS VSS nch l=0.26u w=0.8u
m7690 VSS 3991 VSS VSS nch l=0.26u w=0.8u
m7691 VSS 3992 VSS VSS nch l=0.26u w=0.8u
m7692 VSS 3995 VSS VSS nch l=0.26u w=0.8u
m7693 VSS 3996 VSS VSS nch l=0.26u w=0.8u
m7694 VSS 3999 VSS VSS nch l=0.26u w=0.8u
m7695 VSS 4000 VSS VSS nch l=0.26u w=0.8u
m7696 VSS 4003 VSS VSS nch l=0.26u w=0.8u
m7697 VSS 4004 VSS VSS nch l=0.26u w=0.8u
m7698 VSS 4007 VSS VSS nch l=0.26u w=0.8u
m7699 VSS 4008 VSS VSS nch l=0.26u w=0.8u
m7700 VSS 4011 VSS VSS nch l=0.26u w=0.8u
m7701 VSS 4012 VSS VSS nch l=0.26u w=0.8u
m7702 VSS 4015 VSS VSS nch l=0.26u w=0.8u
m7703 VSS 4016 VSS VSS nch l=0.26u w=0.8u
m7704 VSS 4019 VSS VSS nch l=0.26u w=0.8u
m7705 VSS 4020 VSS VSS nch l=0.26u w=0.8u
m7706 VSS 4023 VSS VSS nch l=0.26u w=0.8u
m7707 VSS 4024 VSS VSS nch l=0.26u w=0.8u
m7708 VSS 4027 VSS VSS nch l=0.26u w=0.8u
m7709 VSS 4028 VSS VSS nch l=0.26u w=0.8u
m7710 VSS 4031 VSS VSS nch l=0.26u w=0.8u
m7711 VSS 4032 VSS VSS nch l=0.26u w=0.8u
m7712 VSS 4035 VSS VSS nch l=0.26u w=0.8u
m7713 VSS 4036 VSS VSS nch l=0.26u w=0.8u
m7714 VSS 4051 71700 VSS nch l=0.04u w=0.12u
m7715 VSS 4328 4046 VSS nch l=0.04u w=0.4u
m7716 VSS 4038 VSS VSS nch l=0.26u w=0.8u
m7717 VSS 4053 4048 VSS nch l=0.04u w=0.4u
m7718 4049 3964 VSS VSS nch l=0.04u w=0.4u
m7719 VSS 4057 4045 VSS nch l=0.04u w=0.4u
m7720 71701 4040 VSS VSS nch l=0.04u w=0.8u
m7721 4051 4041 VSS VSS nch l=0.04u w=0.4u
m7722 CLKSSCG 4047 VSS VSS nch l=0.04u w=0.4u
m7723 71702 3524 VSS VSS nch l=0.04u w=0.8u
m7724 VSS 3971 VSS VSS nch l=0.26u w=0.8u
m7725 VSS 3972 VSS VSS nch l=0.26u w=0.8u
m7726 VSS 3975 VSS VSS nch l=0.26u w=0.8u
m7727 VSS 3976 VSS VSS nch l=0.26u w=0.8u
m7728 VSS 3979 VSS VSS nch l=0.26u w=0.8u
m7729 VSS 3980 VSS VSS nch l=0.26u w=0.8u
m7730 VSS 3983 VSS VSS nch l=0.26u w=0.8u
m7731 VSS 3984 VSS VSS nch l=0.26u w=0.8u
m7732 VSS 3987 VSS VSS nch l=0.26u w=0.8u
m7733 VSS 3988 VSS VSS nch l=0.26u w=0.8u
m7734 VSS 3991 VSS VSS nch l=0.26u w=0.8u
m7735 VSS 3992 VSS VSS nch l=0.26u w=0.8u
m7736 VSS 3995 VSS VSS nch l=0.26u w=0.8u
m7737 VSS 3996 VSS VSS nch l=0.26u w=0.8u
m7738 VSS 3999 VSS VSS nch l=0.26u w=0.8u
m7739 VSS 4000 VSS VSS nch l=0.26u w=0.8u
m7740 VSS 4003 VSS VSS nch l=0.26u w=0.8u
m7741 VSS 4004 VSS VSS nch l=0.26u w=0.8u
m7742 VSS 4007 VSS VSS nch l=0.26u w=0.8u
m7743 VSS 4008 VSS VSS nch l=0.26u w=0.8u
m7744 VSS 4011 VSS VSS nch l=0.26u w=0.8u
m7745 VSS 4012 VSS VSS nch l=0.26u w=0.8u
m7746 VSS 4015 VSS VSS nch l=0.26u w=0.8u
m7747 VSS 4016 VSS VSS nch l=0.26u w=0.8u
m7748 VSS 4019 VSS VSS nch l=0.26u w=0.8u
m7749 VSS 4020 VSS VSS nch l=0.26u w=0.8u
m7750 VSS 4023 VSS VSS nch l=0.26u w=0.8u
m7751 VSS 4024 VSS VSS nch l=0.26u w=0.8u
m7752 VSS 4027 VSS VSS nch l=0.26u w=0.8u
m7753 VSS 4028 VSS VSS nch l=0.26u w=0.8u
m7754 VSS 4031 VSS VSS nch l=0.26u w=0.8u
m7755 VSS 4032 VSS VSS nch l=0.26u w=0.8u
m7756 VSS 4035 VSS VSS nch l=0.26u w=0.8u
m7757 VSS 4036 VSS VSS nch l=0.26u w=0.8u
m7758 VSS 3964 4049 VSS nch l=0.04u w=0.4u
m7759 71703 4045 VSS VSS nch l=0.04u w=0.12u
m7760 71704 3450 71701 VSS nch l=0.04u w=0.8u
m7761 VSS 4038 VSS VSS nch l=0.26u w=0.8u
m7762 4055 4046 3965 VSS nch l=0.04u w=0.4u
m7763 VSS 4047 CLKSSCG VSS nch l=0.04u w=0.4u
m7764 71705 3484 4053 VSS nch l=0.04u w=0.8u
m7765 4054 3959 71702 VSS nch l=0.04u w=0.8u
m7766 4049 3964 VSS VSS nch l=0.04u w=0.4u
m7767 4057 4251 71703 VSS nch l=0.04u w=0.12u
m7768 4050 2969 71704 VSS nch l=0.04u w=0.8u
m7769 4056 4328 4051 VSS nch l=0.04u w=0.4u
m7770 71706 4328 4055 VSS nch l=0.04u w=0.24u
m7771 CLKSSCG 4047 VSS VSS nch l=0.04u w=0.4u
m7772 71707 4351 71705 VSS nch l=0.04u w=0.8u
m7773 71708 3959 4054 VSS nch l=0.04u w=0.8u
m7774 VSS 3971 VSS VSS nch l=0.26u w=0.8u
m7775 VSS 3972 VSS VSS nch l=0.26u w=0.8u
m7776 VSS 3975 VSS VSS nch l=0.26u w=0.8u
m7777 VSS 3976 VSS VSS nch l=0.26u w=0.8u
m7778 VSS 3979 VSS VSS nch l=0.26u w=0.8u
m7779 VSS 3980 VSS VSS nch l=0.26u w=0.8u
m7780 VSS 3983 VSS VSS nch l=0.26u w=0.8u
m7781 VSS 3984 VSS VSS nch l=0.26u w=0.8u
m7782 VSS 3987 VSS VSS nch l=0.26u w=0.8u
m7783 VSS 3988 VSS VSS nch l=0.26u w=0.8u
m7784 VSS 3991 VSS VSS nch l=0.26u w=0.8u
m7785 VSS 3992 VSS VSS nch l=0.26u w=0.8u
m7786 VSS 3995 VSS VSS nch l=0.26u w=0.8u
m7787 VSS 3996 VSS VSS nch l=0.26u w=0.8u
m7788 VSS 3999 VSS VSS nch l=0.26u w=0.8u
m7789 VSS 4000 VSS VSS nch l=0.26u w=0.8u
m7790 VSS 4003 VSS VSS nch l=0.26u w=0.8u
m7791 VSS 4004 VSS VSS nch l=0.26u w=0.8u
m7792 VSS 4007 VSS VSS nch l=0.26u w=0.8u
m7793 VSS 4008 VSS VSS nch l=0.26u w=0.8u
m7794 VSS 4011 VSS VSS nch l=0.26u w=0.8u
m7795 VSS 4012 VSS VSS nch l=0.26u w=0.8u
m7796 VSS 4015 VSS VSS nch l=0.26u w=0.8u
m7797 VSS 4016 VSS VSS nch l=0.26u w=0.8u
m7798 VSS 4019 VSS VSS nch l=0.26u w=0.8u
m7799 VSS 4020 VSS VSS nch l=0.26u w=0.8u
m7800 VSS 4023 VSS VSS nch l=0.26u w=0.8u
m7801 VSS 4024 VSS VSS nch l=0.26u w=0.8u
m7802 VSS 4027 VSS VSS nch l=0.26u w=0.8u
m7803 VSS 4028 VSS VSS nch l=0.26u w=0.8u
m7804 VSS 4031 VSS VSS nch l=0.26u w=0.8u
m7805 VSS 4032 VSS VSS nch l=0.26u w=0.8u
m7806 VSS 4035 VSS VSS nch l=0.26u w=0.8u
m7807 VSS 4036 VSS VSS nch l=0.26u w=0.8u
m7808 VSS 3964 4049 VSS nch l=0.04u w=0.4u
m7809 4058 4059 4057 VSS nch l=0.04u w=0.4u
m7810 VSS 4038 VSS VSS nch l=0.26u w=0.8u
m7811 71709 3966 4056 VSS nch l=0.04u w=0.12u
m7812 VSS 4061 71706 VSS nch l=0.04u w=0.24u
m7813 VSS 4047 CLKSSCG VSS nch l=0.04u w=0.4u
m7814 VSS 4064 71707 VSS nch l=0.04u w=0.8u
m7815 VSS 3524 71708 VSS nch l=0.04u w=0.8u
m7816 4060 4050 VSS VSS nch l=0.04u w=0.4u
m7817 VSS 4063 71709 VSS nch l=0.04u w=0.12u
m7818 71710 4043 VSS VSS nch l=0.04u w=0.8u
m7819 VSS 3971 VSS VSS nch l=0.26u w=0.8u
m7820 VSS 3972 VSS VSS nch l=0.26u w=0.8u
m7821 VSS 3975 VSS VSS nch l=0.26u w=0.8u
m7822 VSS 3976 VSS VSS nch l=0.26u w=0.8u
m7823 VSS 3979 VSS VSS nch l=0.26u w=0.8u
m7824 VSS 3980 VSS VSS nch l=0.26u w=0.8u
m7825 VSS 3983 VSS VSS nch l=0.26u w=0.8u
m7826 VSS 3984 VSS VSS nch l=0.26u w=0.8u
m7827 VSS 3987 VSS VSS nch l=0.26u w=0.8u
m7828 VSS 3988 VSS VSS nch l=0.26u w=0.8u
m7829 VSS 3991 VSS VSS nch l=0.26u w=0.8u
m7830 VSS 3992 VSS VSS nch l=0.26u w=0.8u
m7831 VSS 3995 VSS VSS nch l=0.26u w=0.8u
m7832 VSS 3996 VSS VSS nch l=0.26u w=0.8u
m7833 VSS 3999 VSS VSS nch l=0.26u w=0.8u
m7834 VSS 4000 VSS VSS nch l=0.26u w=0.8u
m7835 VSS 4003 VSS VSS nch l=0.26u w=0.8u
m7836 VSS 4004 VSS VSS nch l=0.26u w=0.8u
m7837 VSS 4007 VSS VSS nch l=0.26u w=0.8u
m7838 VSS 4008 VSS VSS nch l=0.26u w=0.8u
m7839 VSS 4011 VSS VSS nch l=0.26u w=0.8u
m7840 VSS 4012 VSS VSS nch l=0.26u w=0.8u
m7841 VSS 4015 VSS VSS nch l=0.26u w=0.8u
m7842 VSS 4016 VSS VSS nch l=0.26u w=0.8u
m7843 VSS 4019 VSS VSS nch l=0.26u w=0.8u
m7844 VSS 4020 VSS VSS nch l=0.26u w=0.8u
m7845 VSS 4023 VSS VSS nch l=0.26u w=0.8u
m7846 VSS 4024 VSS VSS nch l=0.26u w=0.8u
m7847 VSS 4027 VSS VSS nch l=0.26u w=0.8u
m7848 VSS 4028 VSS VSS nch l=0.26u w=0.8u
m7849 VSS 4031 VSS VSS nch l=0.26u w=0.8u
m7850 VSS 4032 VSS VSS nch l=0.26u w=0.8u
m7851 VSS 4035 VSS VSS nch l=0.26u w=0.8u
m7852 VSS 4036 VSS VSS nch l=0.26u w=0.8u
m7853 4062 4049 VSS VSS nch l=0.04u w=0.4u
m7854 VSS 4038 VSS VSS nch l=0.26u w=0.8u
m7855 VSS 4251 4059 VSS nch l=0.04u w=0.4u
m7856 4063 4056 VSS VSS nch l=0.04u w=0.4u
m7857 4061 4055 71710 VSS nch l=0.04u w=0.8u
m7858 4064 4136 VSS VSS nch l=0.04u w=0.4u
m7859 3117 4054 VSS VSS nch l=0.04u w=0.4u
m7860 VSS 4049 4062 VSS nch l=0.04u w=0.4u
m7861 71713 4060 VSS VSS nch l=0.04u w=0.8u
m7862 VSS 3971 VSS VSS nch l=0.26u w=0.8u
m7863 VSS 3972 VSS VSS nch l=0.26u w=0.8u
m7864 VSS 3975 VSS VSS nch l=0.26u w=0.8u
m7865 VSS 3976 VSS VSS nch l=0.26u w=0.8u
m7866 VSS 3979 VSS VSS nch l=0.26u w=0.8u
m7867 VSS 3980 VSS VSS nch l=0.26u w=0.8u
m7868 VSS 3983 VSS VSS nch l=0.26u w=0.8u
m7869 VSS 3984 VSS VSS nch l=0.26u w=0.8u
m7870 VSS 3987 VSS VSS nch l=0.26u w=0.8u
m7871 VSS 3988 VSS VSS nch l=0.26u w=0.8u
m7872 VSS 3991 VSS VSS nch l=0.26u w=0.8u
m7873 VSS 3992 VSS VSS nch l=0.26u w=0.8u
m7874 VSS 3995 VSS VSS nch l=0.26u w=0.8u
m7875 VSS 3996 VSS VSS nch l=0.26u w=0.8u
m7876 VSS 3999 VSS VSS nch l=0.26u w=0.8u
m7877 VSS 4000 VSS VSS nch l=0.26u w=0.8u
m7878 VSS 4003 VSS VSS nch l=0.26u w=0.8u
m7879 VSS 4004 VSS VSS nch l=0.26u w=0.8u
m7880 VSS 4007 VSS VSS nch l=0.26u w=0.8u
m7881 VSS 4008 VSS VSS nch l=0.26u w=0.8u
m7882 VSS 4011 VSS VSS nch l=0.26u w=0.8u
m7883 VSS 4012 VSS VSS nch l=0.26u w=0.8u
m7884 VSS 4015 VSS VSS nch l=0.26u w=0.8u
m7885 VSS 4016 VSS VSS nch l=0.26u w=0.8u
m7886 VSS 4019 VSS VSS nch l=0.26u w=0.8u
m7887 VSS 4020 VSS VSS nch l=0.26u w=0.8u
m7888 VSS 4023 VSS VSS nch l=0.26u w=0.8u
m7889 VSS 4024 VSS VSS nch l=0.26u w=0.8u
m7890 VSS 4027 VSS VSS nch l=0.26u w=0.8u
m7891 VSS 4028 VSS VSS nch l=0.26u w=0.8u
m7892 VSS 4031 VSS VSS nch l=0.26u w=0.8u
m7893 VSS 4032 VSS VSS nch l=0.26u w=0.8u
m7894 VSS 4035 VSS VSS nch l=0.26u w=0.8u
m7895 VSS 4036 VSS VSS nch l=0.26u w=0.8u
m7896 VSS 4136 4064 VSS nch l=0.04u w=0.4u
m7897 VSS 4038 VSS VSS nch l=0.26u w=0.8u
m7898 4062 4049 VSS VSS nch l=0.04u w=0.4u
m7899 71715 4218 VSS VSS nch l=0.04u w=0.8u
m7900 71716 3484 71713 VSS nch l=0.04u w=0.8u
m7901 4067 4063 VSS VSS nch l=0.04u w=0.4u
m7902 4066 4328 4061 VSS nch l=0.04u w=0.4u
m7903 4068 4069 VSS VSS nch l=0.04u w=0.8u
m7904 4071 4070 VSS VSS nch l=0.04u w=0.8u
m7905 4072 4073 VSS VSS nch l=0.04u w=0.8u
m7906 4075 4074 VSS VSS nch l=0.04u w=0.8u
m7907 4076 4077 VSS VSS nch l=0.04u w=0.8u
m7908 4079 4078 VSS VSS nch l=0.04u w=0.8u
m7909 4080 4081 VSS VSS nch l=0.04u w=0.8u
m7910 4083 4082 VSS VSS nch l=0.04u w=0.8u
m7911 4084 4085 VSS VSS nch l=0.04u w=0.8u
m7912 4087 4086 VSS VSS nch l=0.04u w=0.8u
m7913 4088 4089 VSS VSS nch l=0.04u w=0.8u
m7914 4091 4090 VSS VSS nch l=0.04u w=0.8u
m7915 4092 4093 VSS VSS nch l=0.04u w=0.8u
m7916 4095 4094 VSS VSS nch l=0.04u w=0.8u
m7917 4096 4097 VSS VSS nch l=0.04u w=0.8u
m7918 4099 4098 VSS VSS nch l=0.04u w=0.8u
m7919 4100 4101 VSS VSS nch l=0.04u w=0.8u
m7920 4103 4102 VSS VSS nch l=0.04u w=0.8u
m7921 4104 4105 VSS VSS nch l=0.04u w=0.8u
m7922 4107 4106 VSS VSS nch l=0.04u w=0.8u
m7923 4108 4109 VSS VSS nch l=0.04u w=0.8u
m7924 4111 4110 VSS VSS nch l=0.04u w=0.8u
m7925 4112 4113 VSS VSS nch l=0.04u w=0.8u
m7926 4115 4114 VSS VSS nch l=0.04u w=0.8u
m7927 4116 4117 VSS VSS nch l=0.04u w=0.8u
m7928 4119 4118 VSS VSS nch l=0.04u w=0.8u
m7929 4120 4121 VSS VSS nch l=0.04u w=0.8u
m7930 4123 4122 VSS VSS nch l=0.04u w=0.8u
m7931 4124 4125 VSS VSS nch l=0.04u w=0.8u
m7932 4127 4126 VSS VSS nch l=0.04u w=0.8u
m7933 4128 4129 VSS VSS nch l=0.04u w=0.8u
m7934 4131 4130 VSS VSS nch l=0.04u w=0.8u
m7935 4132 4133 VSS VSS nch l=0.04u w=0.8u
m7936 4135 4134 VSS VSS nch l=0.04u w=0.8u
m7937 71717 4363 VSS VSS nch l=0.04u w=0.8u
m7938 4139 4138 VSS VSS nch l=0.04u w=0.8u
m7939 VSS 4049 4062 VSS nch l=0.04u w=0.4u
m7940 4058 4224 71715 VSS nch l=0.04u w=0.8u
m7941 4065 3953 71716 VSS nch l=0.04u w=0.8u
m7942 71718 4046 4066 VSS nch l=0.04u w=0.12u
m7943 VSS 4216 4136 VSS nch l=0.04u w=0.4u
m7944 4137 4054 71717 VSS nch l=0.04u w=0.8u
m7945 4062 4049 VSS VSS nch l=0.04u w=0.4u
m7946 71719 4224 4058 VSS nch l=0.04u w=0.8u
m7947 VSS 4226 71718 VSS nch l=0.04u w=0.12u
m7948 4212 4230 VSS VSS nch l=0.04u w=0.4u
m7949 VSS 4140 4140 VSS nch l=0.04u w=0.8u
m7950 VSS 4143 4143 VSS nch l=0.04u w=0.8u
m7951 VSS 4144 4144 VSS nch l=0.04u w=0.8u
m7952 VSS 4147 4147 VSS nch l=0.04u w=0.8u
m7953 VSS 4148 4148 VSS nch l=0.04u w=0.8u
m7954 VSS 4151 4151 VSS nch l=0.04u w=0.8u
m7955 VSS 4152 4152 VSS nch l=0.04u w=0.8u
m7956 VSS 4155 4155 VSS nch l=0.04u w=0.8u
m7957 VSS 4156 4156 VSS nch l=0.04u w=0.8u
m7958 VSS 4159 4159 VSS nch l=0.04u w=0.8u
m7959 VSS 4160 4160 VSS nch l=0.04u w=0.8u
m7960 VSS 4163 4163 VSS nch l=0.04u w=0.8u
m7961 VSS 4164 4164 VSS nch l=0.04u w=0.8u
m7962 VSS 4167 4167 VSS nch l=0.04u w=0.8u
m7963 VSS 4168 4168 VSS nch l=0.04u w=0.8u
m7964 VSS 4171 4171 VSS nch l=0.04u w=0.8u
m7965 VSS 4172 4172 VSS nch l=0.04u w=0.8u
m7966 VSS 4175 4175 VSS nch l=0.04u w=0.8u
m7967 VSS 4176 4176 VSS nch l=0.04u w=0.8u
m7968 VSS 4179 4179 VSS nch l=0.04u w=0.8u
m7969 VSS 4180 4180 VSS nch l=0.04u w=0.8u
m7970 VSS 4183 4183 VSS nch l=0.04u w=0.8u
m7971 VSS 4184 4184 VSS nch l=0.04u w=0.8u
m7972 VSS 4187 4187 VSS nch l=0.04u w=0.8u
m7973 VSS 4188 4188 VSS nch l=0.04u w=0.8u
m7974 VSS 4191 4191 VSS nch l=0.04u w=0.8u
m7975 VSS 4192 4192 VSS nch l=0.04u w=0.8u
m7976 VSS 4195 4195 VSS nch l=0.04u w=0.8u
m7977 VSS 4196 4196 VSS nch l=0.04u w=0.8u
m7978 VSS 4199 4199 VSS nch l=0.04u w=0.8u
m7979 VSS 4200 4200 VSS nch l=0.04u w=0.8u
m7980 VSS 4203 4203 VSS nch l=0.04u w=0.8u
m7981 VSS 4204 4204 VSS nch l=0.04u w=0.8u
m7982 VSS 4207 4207 VSS nch l=0.04u w=0.8u
m7983 VSS 4208 4208 VSS nch l=0.04u w=0.8u
m7984 71720 4136 VSS VSS nch l=0.04u w=0.12u
m7985 VSS 4049 4062 VSS nch l=0.04u w=0.4u
m7986 VSS 4211 4211 VSS nch l=0.04u w=0.8u
m7987 VSS 4218 71719 VSS nch l=0.04u w=0.8u
m7988 4213 4065 VSS VSS nch l=0.04u w=0.4u
m7989 4214 4066 VSS VSS nch l=0.04u w=0.4u
m7990 4216 4234 71720 VSS nch l=0.04u w=0.12u
m7991 4217 4617 VSS VSS nch l=0.04u w=0.4u
m7992 VSS 4328 4215 VSS nch l=0.04u w=0.4u
m7993 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m7994 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m7995 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m7996 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m7997 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m7998 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m7999 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8000 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8001 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8002 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8003 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8004 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8005 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8006 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8007 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8008 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8009 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8010 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8011 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8012 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8013 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8014 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8015 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8016 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8017 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8018 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8019 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8020 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8021 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8022 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8023 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8024 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8025 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8026 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8027 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8028 4220 4251 4216 VSS nch l=0.04u w=0.4u
m8029 VSS 4210 VSS VSS nch l=0.26u w=0.8u
m8030 4062 4049 VSS VSS nch l=0.04u w=0.4u
m8031 71721 4238 4218 VSS nch l=0.04u w=0.8u
m8032 4219 4221 4065 VSS nch l=0.04u w=0.4u
m8033 71722 4043 VSS VSS nch l=0.04u w=0.8u
m8034 4222 4217 4137 VSS nch l=0.04u w=0.4u
m8035 VSS 4049 4062 VSS nch l=0.04u w=0.4u
m8036 VSS 4232 71721 VSS nch l=0.04u w=0.8u
m8037 4221 4065 4219 VSS nch l=0.04u w=0.4u
m8038 69 4214 71722 VSS nch l=0.04u w=0.8u
m8039 4223 4215 4067 VSS nch l=0.04u w=0.4u
m8040 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m8041 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m8042 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m8043 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m8044 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m8045 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m8046 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8047 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8048 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8049 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8050 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8051 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8052 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8053 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8054 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8055 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8056 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8057 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8058 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8059 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8060 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8061 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8062 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8063 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8064 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8065 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8066 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8067 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8068 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8069 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8070 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8071 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8072 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8073 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8074 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8075 VSS 4210 VSS VSS nch l=0.26u w=0.8u
m8076 VSS 4227 4220 VSS nch l=0.04u w=0.4u
m8077 71723 4617 4222 VSS nch l=0.04u w=0.12u
m8078 4062 4049 VSS VSS nch l=0.04u w=0.4u
m8079 71724 4328 4223 VSS nch l=0.04u w=0.24u
m8080 71725 4220 VSS VSS nch l=0.04u w=0.12u
m8081 VSS 4228 71723 VSS nch l=0.04u w=0.12u
m8082 VSS 4049 4062 VSS nch l=0.04u w=0.4u
m8083 71726 911 4224 VSS nch l=0.04u w=0.8u
m8084 4225 4062 VSS VSS nch l=0.04u w=0.4u
m8085 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m8086 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m8087 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m8088 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m8089 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m8090 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m8091 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8092 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8093 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8094 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8095 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8096 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8097 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8098 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8099 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8100 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8101 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8102 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8103 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8104 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8105 4226 69 VSS VSS nch l=0.04u w=0.4u
m8106 VSS 4229 71724 VSS nch l=0.04u w=0.24u
m8107 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8108 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8109 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8110 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8111 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8112 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8113 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8114 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8115 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8116 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8117 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8118 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8119 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8120 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8121 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8122 VSS 4210 VSS VSS nch l=0.26u w=0.8u
m8123 4227 4251 71725 VSS nch l=0.04u w=0.12u
m8124 4228 4222 VSS VSS nch l=0.04u w=0.4u
m8125 4062 4049 VSS VSS nch l=0.04u w=0.4u
m8126 VSS 4062 71726 VSS nch l=0.04u w=0.8u
m8127 71727 4212 VSS VSS nch l=0.04u w=0.8u
m8128 4231 4234 4227 VSS nch l=0.04u w=0.4u
m8129 VSS 4049 4062 VSS nch l=0.04u w=0.4u
m8130 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m8131 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m8132 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m8133 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m8134 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m8135 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m8136 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8137 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8138 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8139 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8140 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8141 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8142 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8143 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8144 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8145 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8146 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8147 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8148 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8149 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8150 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8151 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8152 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8153 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8154 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8155 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8156 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8157 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8158 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8159 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8160 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8161 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8162 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8163 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8164 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8165 4229 4223 71727 VSS nch l=0.04u w=0.8u
m8166 71728 4062 VSS VSS nch l=0.04u w=0.8u
m8167 VSS 2616 4230 VSS nch l=0.04u w=0.4u
m8168 VSS 4210 VSS VSS nch l=0.26u w=0.8u
m8169 4235 4617 4228 VSS nch l=0.04u w=0.4u
m8170 VSS 4062 4232 VSS nch l=0.04u w=0.4u
m8171 4233 2501 71728 VSS nch l=0.04u w=0.8u
m8172 VSS 4251 4234 VSS nch l=0.04u w=0.4u
m8173 71730 4217 4235 VSS nch l=0.04u w=0.12u
m8174 4236 4251 VSS VSS nch l=0.04u w=0.4u
m8175 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m8176 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m8177 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m8178 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m8179 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m8180 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m8181 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8182 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8183 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8184 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8185 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8186 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8187 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8188 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8189 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8190 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8191 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8192 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8193 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8194 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8195 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8196 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8197 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8198 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8199 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8200 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8201 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8202 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8203 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8204 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8205 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8206 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8207 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8208 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8209 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8210 4237 4328 4229 VSS nch l=0.04u w=0.4u
m8211 VSS 4210 VSS VSS nch l=0.26u w=0.8u
m8212 VSS 4242 71730 VSS nch l=0.04u w=0.12u
m8213 4238 PD 3963 VSS nch l=0.04u w=0.4u
m8214 71732 4215 4237 VSS nch l=0.04u w=0.12u
m8215 71733 4225 VSS VSS nch l=0.04u w=0.8u
m8216 4241 4240 VSS VSS nch l=0.04u w=0.8u
m8217 71735 4250 VSS VSS nch l=0.04u w=0.8u
m8218 4242 4235 VSS VSS nch l=0.04u w=0.4u
m8219 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m8220 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m8221 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m8222 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m8223 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m8224 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m8225 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8226 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8227 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8228 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8229 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8230 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8231 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8232 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8233 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8234 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8235 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8236 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8237 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8238 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8239 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8240 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8241 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8242 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8243 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8244 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8245 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8246 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8247 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8248 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8249 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8250 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8251 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8252 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8253 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8254 4243 4236 4062 VSS nch l=0.04u w=0.4u
m8255 PD 3963 4238 VSS nch l=0.04u w=0.4u
m8256 VSS 4324 71732 VSS nch l=0.04u w=0.12u
m8257 4239 4219 71733 VSS nch l=0.04u w=0.8u
m8258 4231 4325 71735 VSS nch l=0.04u w=0.8u
m8259 71737 4251 4243 VSS nch l=0.04u w=0.12u
m8260 4244 4237 VSS VSS nch l=0.04u w=0.4u
m8261 71739 4325 4231 VSS nch l=0.04u w=0.8u
m8262 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m8263 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m8264 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m8265 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m8266 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m8267 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m8268 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8269 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8270 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8271 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8272 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8273 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8274 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8275 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8276 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8277 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8278 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8279 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8280 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8281 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8282 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8283 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8284 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8285 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8286 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8287 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8288 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8289 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8290 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8291 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8292 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8293 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8294 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8295 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8296 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8297 71740 4242 VSS VSS nch l=0.04u w=0.8u
m8298 VSS 4249 71737 VSS nch l=0.04u w=0.12u
m8299 VSS PD 4245 VSS nch l=0.04u w=0.4u
m8300 71741 4239 VSS VSS nch l=0.04u w=0.8u
m8301 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8302 VSS 4250 71739 VSS nch l=0.04u w=0.8u
m8303 4246 4359 71740 VSS nch l=0.04u w=0.8u
m8304 4249 4243 VSS VSS nch l=0.04u w=0.4u
m8305 71743 4212 VSS VSS nch l=0.04u w=0.8u
m8306 4247 4233 71741 VSS nch l=0.04u w=0.8u
m8307 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8308 VSS 4141 VSS VSS nch l=0.26u w=0.8u
m8309 VSS 4142 VSS VSS nch l=0.26u w=0.8u
m8310 VSS 4145 VSS VSS nch l=0.26u w=0.8u
m8311 VSS 4146 VSS VSS nch l=0.26u w=0.8u
m8312 VSS 4149 VSS VSS nch l=0.26u w=0.8u
m8313 VSS 4150 VSS VSS nch l=0.26u w=0.8u
m8314 VSS 4153 VSS VSS nch l=0.26u w=0.8u
m8315 VSS 4154 VSS VSS nch l=0.26u w=0.8u
m8316 VSS 4157 VSS VSS nch l=0.26u w=0.8u
m8317 VSS 4158 VSS VSS nch l=0.26u w=0.8u
m8318 VSS 4161 VSS VSS nch l=0.26u w=0.8u
m8319 VSS 4162 VSS VSS nch l=0.26u w=0.8u
m8320 VSS 4165 VSS VSS nch l=0.26u w=0.8u
m8321 VSS 4166 VSS VSS nch l=0.26u w=0.8u
m8322 VSS 4169 VSS VSS nch l=0.26u w=0.8u
m8323 VSS 4170 VSS VSS nch l=0.26u w=0.8u
m8324 VSS 4173 VSS VSS nch l=0.26u w=0.8u
m8325 VSS 4174 VSS VSS nch l=0.26u w=0.8u
m8326 VSS 4177 VSS VSS nch l=0.26u w=0.8u
m8327 VSS 4178 VSS VSS nch l=0.26u w=0.8u
m8328 VSS 4181 VSS VSS nch l=0.26u w=0.8u
m8329 VSS 4182 VSS VSS nch l=0.26u w=0.8u
m8330 VSS 4185 VSS VSS nch l=0.26u w=0.8u
m8331 VSS 4186 VSS VSS nch l=0.26u w=0.8u
m8332 VSS 4189 VSS VSS nch l=0.26u w=0.8u
m8333 VSS 4190 VSS VSS nch l=0.26u w=0.8u
m8334 VSS 4193 VSS VSS nch l=0.26u w=0.8u
m8335 VSS 4194 VSS VSS nch l=0.26u w=0.8u
m8336 VSS 4197 VSS VSS nch l=0.26u w=0.8u
m8337 VSS 4198 VSS VSS nch l=0.26u w=0.8u
m8338 VSS 4201 VSS VSS nch l=0.26u w=0.8u
m8339 VSS 4202 VSS VSS nch l=0.26u w=0.8u
m8340 VSS 4205 VSS VSS nch l=0.26u w=0.8u
m8341 VSS 4206 VSS VSS nch l=0.26u w=0.8u
m8342 VSS 4209 VSS VSS nch l=0.26u w=0.8u
m8343 70 4244 71743 VSS nch l=0.04u w=0.8u
m8344 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8345 71745 4233 4247 VSS nch l=0.04u w=0.8u
m8346 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8347 4252 4253 VSS VSS nch l=0.04u w=0.8u
m8348 4255 4254 VSS VSS nch l=0.04u w=0.8u
m8349 4256 4257 VSS VSS nch l=0.04u w=0.8u
m8350 4259 4258 VSS VSS nch l=0.04u w=0.8u
m8351 4260 4261 VSS VSS nch l=0.04u w=0.8u
m8352 4263 4262 VSS VSS nch l=0.04u w=0.8u
m8353 4264 4265 VSS VSS nch l=0.04u w=0.8u
m8354 4267 4266 VSS VSS nch l=0.04u w=0.8u
m8355 4268 4269 VSS VSS nch l=0.04u w=0.8u
m8356 4271 4270 VSS VSS nch l=0.04u w=0.8u
m8357 4272 4273 VSS VSS nch l=0.04u w=0.8u
m8358 4275 4274 VSS VSS nch l=0.04u w=0.8u
m8359 4276 4277 VSS VSS nch l=0.04u w=0.8u
m8360 4279 4278 VSS VSS nch l=0.04u w=0.8u
m8361 4280 4281 VSS VSS nch l=0.04u w=0.8u
m8362 4283 4282 VSS VSS nch l=0.04u w=0.8u
m8363 4284 4285 VSS VSS nch l=0.04u w=0.8u
m8364 4287 4286 VSS VSS nch l=0.04u w=0.8u
m8365 4288 4289 VSS VSS nch l=0.04u w=0.8u
m8366 4291 4290 VSS VSS nch l=0.04u w=0.8u
m8367 4292 4293 VSS VSS nch l=0.04u w=0.8u
m8368 4295 4294 VSS VSS nch l=0.04u w=0.8u
m8369 4296 4297 VSS VSS nch l=0.04u w=0.8u
m8370 4299 4298 VSS VSS nch l=0.04u w=0.8u
m8371 4300 4301 VSS VSS nch l=0.04u w=0.8u
m8372 4303 4302 VSS VSS nch l=0.04u w=0.8u
m8373 4304 4305 VSS VSS nch l=0.04u w=0.8u
m8374 4307 4306 VSS VSS nch l=0.04u w=0.8u
m8375 4308 4309 VSS VSS nch l=0.04u w=0.8u
m8376 4311 4310 VSS VSS nch l=0.04u w=0.8u
m8377 4312 4313 VSS VSS nch l=0.04u w=0.8u
m8378 4315 4314 VSS VSS nch l=0.04u w=0.8u
m8379 4316 4317 VSS VSS nch l=0.04u w=0.8u
m8380 4319 4318 VSS VSS nch l=0.04u w=0.8u
m8381 4320 4321 VSS VSS nch l=0.04u w=0.8u
m8382 71747 4337 4250 VSS nch l=0.04u w=0.8u
m8383 4322 4617 VSS VSS nch l=0.04u w=0.4u
m8384 4323 4249 VSS VSS nch l=0.04u w=0.4u
m8385 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8386 VSS 4239 71745 VSS nch l=0.04u w=0.8u
m8387 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8388 VSS 4331 71747 VSS nch l=0.04u w=0.8u
m8389 VSS 4249 4323 VSS nch l=0.04u w=0.4u
m8390 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8391 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8392 4324 70 VSS VSS nch l=0.04u w=0.4u
m8393 4326 4322 4246 VSS nch l=0.04u w=0.4u
m8394 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8395 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8396 4327 4251 VSS VSS nch l=0.04u w=0.4u
m8397 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8398 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8399 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8400 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8401 71786 2952 4325 VSS nch l=0.04u w=0.8u
m8402 71787 4617 4326 VSS nch l=0.04u w=0.12u
m8403 4329 4062 VSS VSS nch l=0.04u w=0.4u
m8404 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8405 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8406 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8407 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8408 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8409 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8410 VSS 4062 71786 VSS nch l=0.04u w=0.8u
m8411 VSS 4332 71787 VSS nch l=0.04u w=0.12u
m8412 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8413 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8414 4330 4327 4247 VSS nch l=0.04u w=0.4u
m8415 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8416 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8417 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8418 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8419 4332 4326 VSS VSS nch l=0.04u w=0.4u
m8420 4333 4251 VSS VSS nch l=0.04u w=0.4u
m8421 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8422 71824 4251 4330 VSS nch l=0.04u w=0.12u
m8423 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8424 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8425 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8426 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8427 VSS 4062 4331 VSS nch l=0.04u w=0.4u
m8428 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8429 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8430 VSS 4336 71824 VSS nch l=0.04u w=0.12u
m8431 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8432 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8433 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8434 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8435 4334 4617 4332 VSS nch l=0.04u w=0.4u
m8436 4335 4333 4329 VSS nch l=0.04u w=0.4u
m8437 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8438 4336 4330 VSS VSS nch l=0.04u w=0.4u
m8439 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8440 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8441 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8442 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8443 4337 4338 4136 VSS nch l=0.04u w=0.4u
m8444 71825 4322 4334 VSS nch l=0.04u w=0.12u
m8445 71826 4251 4335 VSS nch l=0.04u w=0.12u
m8446 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8447 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8448 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8449 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8450 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8451 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8452 4338 4136 4337 VSS nch l=0.04u w=0.4u
m8453 VSS 4340 71825 VSS nch l=0.04u w=0.12u
m8454 VSS 4342 71826 VSS nch l=0.04u w=0.12u
m8455 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8456 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8457 4339 4251 4336 VSS nch l=0.04u w=0.4u
m8458 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8459 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8460 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8461 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8462 4340 4334 VSS VSS nch l=0.04u w=0.4u
m8463 4342 4335 VSS VSS nch l=0.04u w=0.4u
m8464 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8465 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8466 71827 4327 4339 VSS nch l=0.04u w=0.12u
m8467 VSS 4338 4341 VSS nch l=0.04u w=0.4u
m8468 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8469 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8470 VSS 4221 71827 VSS nch l=0.04u w=0.12u
m8471 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8472 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8473 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8474 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8475 4343 4617 VSS VSS nch l=0.04u w=0.4u
m8476 4344 4251 4342 VSS nch l=0.04u w=0.4u
m8477 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8478 4248 4346 VSS VSS nch l=0.04u w=0.4u
m8479 4221 4339 VSS VSS nch l=0.04u w=0.4u
m8480 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8481 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8482 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8483 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8484 71828 3953 4338 VSS nch l=0.04u w=0.8u
m8485 71829 4333 4344 VSS nch l=0.04u w=0.12u
m8486 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8487 VSS 4346 4248 VSS nch l=0.04u w=0.4u
m8488 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8489 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8490 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8491 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8492 71830 3484 71828 VSS nch l=0.04u w=0.8u
m8493 4345 4343 4340 VSS nch l=0.04u w=0.4u
m8494 VSS 4348 71829 VSS nch l=0.04u w=0.12u
m8495 4251 4362 VSS VSS nch l=0.04u w=0.4u
m8496 4347 4221 VSS VSS nch l=0.04u w=0.4u
m8497 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8498 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8499 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8500 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8501 VSS 4351 71830 VSS nch l=0.04u w=0.8u
m8502 71831 4617 4345 VSS nch l=0.04u w=0.12u
m8503 4348 4344 VSS VSS nch l=0.04u w=0.4u
m8504 VSS 4362 4251 VSS nch l=0.04u w=0.4u
m8505 4349 4368 4346 VSS nch l=0.04u w=0.8u
m8506 VSS 4221 4347 VSS nch l=0.04u w=0.4u
m8507 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8508 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8509 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8510 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8511 VSS 4350 71831 VSS nch l=0.04u w=0.12u
m8512 4346 4368 4349 VSS nch l=0.04u w=0.8u
m8513 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8514 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8515 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8516 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8517 4350 4345 VSS VSS nch l=0.04u w=0.4u
m8518 4351 4357 VSS VSS nch l=0.04u w=0.4u
m8519 4352 4251 VSS VSS nch l=0.04u w=0.4u
m8520 4353 4362 VSS VSS nch l=0.04u w=0.4u
m8521 4349 4368 4346 VSS nch l=0.04u w=0.8u
m8522 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8523 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8524 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8525 4328 4248 VSS VSS nch l=0.04u w=0.4u
m8526 VSS 4357 4351 VSS nch l=0.04u w=0.4u
m8527 VSS 4362 4353 VSS nch l=0.04u w=0.4u
m8528 VSS 4367 4349 VSS nch l=0.04u w=0.8u
m8529 VSS 4354 4354 VSS nch l=0.04u w=0.8u
m8530 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8531 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8532 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8533 VSS 4248 4328 VSS nch l=0.04u w=0.4u
m8534 4356 4617 4350 VSS nch l=0.04u w=0.4u
m8535 4353 4362 VSS VSS nch l=0.04u w=0.4u
m8536 4358 4352 4348 VSS nch l=0.04u w=0.4u
m8537 4349 4367 VSS VSS nch l=0.04u w=0.8u
m8538 71838 4343 4356 VSS nch l=0.04u w=0.12u
m8539 71839 2969 4357 VSS nch l=0.04u w=0.8u
m8540 VSS 4362 4353 VSS nch l=0.04u w=0.4u
m8541 71840 4251 4358 VSS nch l=0.04u w=0.12u
m8542 VSS 4367 4349 VSS nch l=0.04u w=0.8u
m8543 VSS 4355 VSS VSS nch l=0.26u w=0.8u
m8544 VSS 4359 71838 VSS nch l=0.04u w=0.12u
m8545 VSS 4360 71839 VSS nch l=0.04u w=0.8u
m8546 VSS 4361 71840 VSS nch l=0.04u w=0.12u
m8547 4349 4367 VSS VSS nch l=0.04u w=0.8u
m8548 4359 4356 VSS VSS nch l=0.04u w=0.4u
m8549 4361 4358 VSS VSS nch l=0.04u w=0.4u
m8550 VSS 4367 4349 VSS nch l=0.04u w=0.8u
m8551 4362 4366 VSS VSS nch l=0.04u w=0.4u
m8552 VSS 4355 VSS VSS nch l=0.26u w=0.8u
m8553 VSS 4365 4360 VSS nch l=0.04u w=0.4u
m8554 4349 4367 VSS VSS nch l=0.04u w=0.8u
m8555 VSS 4366 4362 VSS nch l=0.04u w=0.4u
m8556 4363 4359 VSS VSS nch l=0.04u w=0.4u
m8557 VSS 4367 4349 VSS nch l=0.04u w=0.8u
m8558 4362 4366 VSS VSS nch l=0.04u w=0.4u
m8559 VSS 4355 VSS VSS nch l=0.26u w=0.8u
m8560 4364 4251 4361 VSS nch l=0.04u w=0.4u
m8561 4349 4367 VSS VSS nch l=0.04u w=0.8u
m8562 VSS 4366 4362 VSS nch l=0.04u w=0.4u
m8563 71859 3450 4365 VSS nch l=0.04u w=0.8u
m8564 71860 4352 4364 VSS nch l=0.04u w=0.12u
m8565 VSS 4355 VSS VSS nch l=0.26u w=0.8u
m8566 4366 4363 VSS VSS nch l=0.04u w=0.4u
m8567 4362 4366 VSS VSS nch l=0.04u w=0.4u
m8568 71865 4040 71859 VSS nch l=0.04u w=0.8u
m8569 VSS 4368 71860 VSS nch l=0.04u w=0.12u
m8570 VSS 4363 4366 VSS nch l=0.04u w=0.4u
m8571 VSS 4366 4362 VSS nch l=0.04u w=0.4u
m8572 VSS 4347 71865 VSS nch l=0.04u w=0.8u
m8573 4368 4364 VSS VSS nch l=0.04u w=0.4u
m8574 VSS DSMPD 4367 VSS nch l=0.04u w=0.4u
m8575 VSS 4355 VSS VSS nch l=0.26u w=0.8u
m8576 4369 4370 VSS VSS nch l=0.04u w=0.8u
m8577 VSS 4372 4372 VSS nch l=0.04u w=0.8u
m8578 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8579 VSS 4374 4374 VSS nch l=0.04u w=0.8u
m8580 VSS 4377 4377 VSS nch l=0.04u w=0.8u
m8581 VSS 4378 4378 VSS nch l=0.04u w=0.8u
m8582 VSS 4381 4381 VSS nch l=0.04u w=0.8u
m8583 VSS 4382 4382 VSS nch l=0.04u w=0.8u
m8584 VSS 4385 4385 VSS nch l=0.04u w=0.8u
m8585 VSS 4386 4386 VSS nch l=0.04u w=0.8u
m8586 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8587 4388 2427 VSS VSS nch l=0.04u w=0.4u
m8588 4389 4390 VSS VSS nch l=0.04u w=0.8u
m8589 VSS 2427 4388 VSS nch l=0.04u w=0.4u
m8590 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8591 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8592 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8593 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8594 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8595 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8596 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8597 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8598 4391 FBDIV[10] VSS VSS nch l=0.04u w=0.4u
m8599 4392 2426 VSS VSS nch l=0.04u w=0.4u
m8600 VSS FBDIV[11] 4391 VSS nch l=0.04u w=0.4u
m8601 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8602 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8603 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8604 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8605 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8606 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8607 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8608 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8609 VSS 2426 4392 VSS nch l=0.04u w=0.4u
m8610 4393 2952 VSS VSS nch l=0.04u w=0.4u
m8611 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8612 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8613 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8614 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8615 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8616 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8617 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8618 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8619 4394 4323 VSS VSS nch l=0.04u w=0.4u
m8620 VSS FBDIV[9] 4393 VSS nch l=0.04u w=0.4u
m8621 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8622 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8623 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8624 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8625 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8626 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8627 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8628 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8629 4395 4394 VSS VSS nch l=0.04u w=0.4u
m8630 71922 4393 VSS VSS nch l=0.04u w=0.8u
m8631 VSS 4394 4395 VSS nch l=0.04u w=0.4u
m8632 4396 4391 71922 VSS nch l=0.04u w=0.8u
m8633 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8634 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8635 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8636 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8637 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8638 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8639 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8640 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8641 4395 4394 VSS VSS nch l=0.04u w=0.4u
m8642 VSS 4394 4395 VSS nch l=0.04u w=0.4u
m8643 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8644 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8645 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8646 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8647 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8648 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8649 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8650 4397 2427 VSS VSS nch l=0.04u w=0.4u
m8651 VSS 4371 VSS VSS nch l=0.26u w=0.8u
m8652 4399 4398 VSS VSS nch l=0.04u w=0.8u
m8653 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8654 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8655 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8656 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8657 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8658 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8659 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8660 4400 3293 VSS VSS nch l=0.04u w=0.4u
m8661 71923 DSMPD VSS VSS nch l=0.04u w=0.8u
m8662 VSS 3783 4400 VSS nch l=0.04u w=0.4u
m8663 71924 4396 71923 VSS nch l=0.04u w=0.8u
m8664 VSS 4403 4403 VSS nch l=0.04u w=0.8u
m8665 VSS 4375 VSS VSS nch l=0.26u w=0.8u
m8666 VSS 4376 VSS VSS nch l=0.26u w=0.8u
m8667 VSS 4379 VSS VSS nch l=0.26u w=0.8u
m8668 VSS 4380 VSS VSS nch l=0.26u w=0.8u
m8669 VSS 4383 VSS VSS nch l=0.26u w=0.8u
m8670 VSS 4384 VSS VSS nch l=0.26u w=0.8u
m8671 VSS 4387 VSS VSS nch l=0.26u w=0.8u
m8672 4401 4397 71924 VSS nch l=0.04u w=0.8u
m8673 4404 4405 VSS VSS nch l=0.04u w=0.8u
m8674 4407 4406 VSS VSS nch l=0.04u w=0.8u
m8675 4408 4409 VSS VSS nch l=0.04u w=0.8u
m8676 4411 4410 VSS VSS nch l=0.04u w=0.8u
m8677 4412 4413 VSS VSS nch l=0.04u w=0.8u
m8678 4415 4414 VSS VSS nch l=0.04u w=0.8u
m8679 4416 4417 VSS VSS nch l=0.04u w=0.8u
m8680 4418 4400 VSS VSS nch l=0.04u w=0.4u
m8681 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8682 71930 DSMPD VSS VSS nch l=0.04u w=0.8u
m8683 VSS 4419 4419 VSS nch l=0.04u w=0.8u
m8684 VSS 4422 4422 VSS nch l=0.04u w=0.8u
m8685 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8686 4424 3480 VSS VSS nch l=0.04u w=0.4u
m8687 71931 4396 71930 VSS nch l=0.04u w=0.8u
m8688 VSS 3937 4424 VSS nch l=0.04u w=0.4u
m8689 4423 2426 71931 VSS nch l=0.04u w=0.8u
m8690 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8691 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8692 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8693 4425 4424 VSS VSS nch l=0.04u w=0.4u
m8694 4426 4423 VSS VSS nch l=0.04u w=0.4u
m8695 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8696 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8697 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8698 71939 4395 VSS VSS nch l=0.04u w=0.8u
m8699 71940 4395 VSS VSS nch l=0.04u w=0.8u
m8700 71941 4395 VSS VSS nch l=0.04u w=0.8u
m8701 71942 4395 VSS VSS nch l=0.04u w=0.8u
m8702 71943 4395 VSS VSS nch l=0.04u w=0.8u
m8703 4432 4467 VSS VSS nch l=0.04u w=0.4u
m8704 4433 4468 VSS VSS nch l=0.04u w=0.4u
m8705 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8706 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8707 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8708 4427 2509 71939 VSS nch l=0.04u w=0.8u
m8709 4428 2747 71940 VSS nch l=0.04u w=0.8u
m8710 4429 3019 71941 VSS nch l=0.04u w=0.8u
m8711 4430 4418 71942 VSS nch l=0.04u w=0.8u
m8712 4431 3783 71943 VSS nch l=0.04u w=0.8u
m8713 VSS 4467 4432 VSS nch l=0.04u w=0.4u
m8714 VSS 4468 4433 VSS nch l=0.04u w=0.4u
m8715 4432 4467 VSS VSS nch l=0.04u w=0.4u
m8716 4433 4468 VSS VSS nch l=0.04u w=0.4u
m8717 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8718 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8719 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8720 VSS 4467 4432 VSS nch l=0.04u w=0.4u
m8721 VSS 4468 4433 VSS nch l=0.04u w=0.4u
m8722 4434 DACPD VSS VSS nch l=0.04u w=0.4u
m8723 4435 DACPD VSS VSS nch l=0.04u w=0.4u
m8724 4436 DACPD VSS VSS nch l=0.04u w=0.4u
m8725 4437 DACPD VSS VSS nch l=0.04u w=0.4u
m8726 4438 DACPD VSS VSS nch l=0.04u w=0.4u
m8727 4432 4467 VSS VSS nch l=0.04u w=0.4u
m8728 4433 4468 VSS VSS nch l=0.04u w=0.4u
m8729 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8730 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8731 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8732 VSS 4467 4432 VSS nch l=0.04u w=0.4u
m8733 VSS 4468 4433 VSS nch l=0.04u w=0.4u
m8734 71944 DACPD VSS VSS nch l=0.04u w=0.8u
m8735 71945 DACPD VSS VSS nch l=0.04u w=0.8u
m8736 71946 DACPD VSS VSS nch l=0.04u w=0.8u
m8737 71947 DACPD VSS VSS nch l=0.04u w=0.8u
m8738 71948 DACPD VSS VSS nch l=0.04u w=0.8u
m8739 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8740 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8741 4439 DACPD 71944 VSS nch l=0.04u w=0.8u
m8742 4440 DACPD 71945 VSS nch l=0.04u w=0.8u
m8743 4441 DACPD 71946 VSS nch l=0.04u w=0.8u
m8744 4442 DACPD 71947 VSS nch l=0.04u w=0.8u
m8745 4443 DACPD 71948 VSS nch l=0.04u w=0.8u
m8746 VSS 4402 VSS VSS nch l=0.26u w=0.8u
m8747 4432 4467 VSS VSS nch l=0.04u w=0.4u
m8748 4433 4468 VSS VSS nch l=0.04u w=0.4u
m8749 4446 4445 VSS VSS nch l=0.04u w=0.8u
m8750 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8751 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8752 VSS 4467 4432 VSS nch l=0.04u w=0.4u
m8753 VSS 4468 4433 VSS nch l=0.04u w=0.4u
m8754 71949 4434 VSS VSS nch l=0.04u w=0.8u
m8755 71950 4435 VSS VSS nch l=0.04u w=0.8u
m8756 71951 4436 VSS VSS nch l=0.04u w=0.8u
m8757 71952 4437 VSS VSS nch l=0.04u w=0.8u
m8758 71953 4438 VSS VSS nch l=0.04u w=0.8u
m8759 4432 4467 VSS VSS nch l=0.04u w=0.4u
m8760 4433 4468 VSS VSS nch l=0.04u w=0.4u
m8761 4447 4427 71949 VSS nch l=0.04u w=0.8u
m8762 4448 4428 71950 VSS nch l=0.04u w=0.8u
m8763 4449 4429 71951 VSS nch l=0.04u w=0.8u
m8764 4450 4430 71952 VSS nch l=0.04u w=0.8u
m8765 4451 4431 71953 VSS nch l=0.04u w=0.8u
m8766 VSS 4453 4453 VSS nch l=0.04u w=0.8u
m8767 VSS 4420 VSS VSS nch l=0.26u w=0.8u
m8768 VSS 4421 VSS VSS nch l=0.26u w=0.8u
m8769 VSS 4467 4432 VSS nch l=0.04u w=0.4u
m8770 VSS 4468 4433 VSS nch l=0.04u w=0.4u
m8771 4454 4455 VSS VSS nch l=0.04u w=0.8u
m8772 4457 4456 VSS VSS nch l=0.04u w=0.8u
m8773 4432 4467 VSS VSS nch l=0.04u w=0.4u
m8774 4433 4468 VSS VSS nch l=0.04u w=0.4u
m8775 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8776 71954 4447 VSS VSS nch l=0.04u w=0.8u
m8777 71955 4448 VSS VSS nch l=0.04u w=0.8u
m8778 71956 4449 VSS VSS nch l=0.04u w=0.8u
m8779 71957 4450 VSS VSS nch l=0.04u w=0.8u
m8780 71958 4451 VSS VSS nch l=0.04u w=0.8u
m8781 VSS 4467 4432 VSS nch l=0.04u w=0.4u
m8782 VSS 4468 4433 VSS nch l=0.04u w=0.4u
m8783 4458 4439 71954 VSS nch l=0.04u w=0.8u
m8784 4459 4440 71955 VSS nch l=0.04u w=0.8u
m8785 4460 4441 71956 VSS nch l=0.04u w=0.8u
m8786 4461 4442 71957 VSS nch l=0.04u w=0.8u
m8787 4462 4443 71958 VSS nch l=0.04u w=0.8u
m8788 VSS 4463 4463 VSS nch l=0.04u w=0.8u
m8789 VSS 4466 4466 VSS nch l=0.04u w=0.8u
m8790 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8791 4467 4480 VSS VSS nch l=0.04u w=0.4u
m8792 4468 4481 VSS VSS nch l=0.04u w=0.4u
m8793 4469 155 VSS VSS nch l=0.04u w=0.4u
m8794 4470 155 VSS VSS nch l=0.04u w=0.4u
m8795 4471 155 VSS VSS nch l=0.04u w=0.4u
m8796 4472 155 VSS VSS nch l=0.04u w=0.4u
m8797 4473 155 VSS VSS nch l=0.04u w=0.4u
m8798 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8799 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8800 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8801 VSS 4480 4467 VSS nch l=0.04u w=0.4u
m8802 VSS 4481 4468 VSS nch l=0.04u w=0.4u
m8803 4467 4480 VSS VSS nch l=0.04u w=0.4u
m8804 4468 4481 VSS VSS nch l=0.04u w=0.4u
m8805 71959 155 VSS VSS nch l=0.04u w=0.8u
m8806 71960 155 VSS VSS nch l=0.04u w=0.8u
m8807 71961 155 VSS VSS nch l=0.04u w=0.8u
m8808 71962 155 VSS VSS nch l=0.04u w=0.8u
m8809 71963 155 VSS VSS nch l=0.04u w=0.8u
m8810 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8811 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8812 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8813 VSS 4480 4467 VSS nch l=0.04u w=0.4u
m8814 VSS 4481 4468 VSS nch l=0.04u w=0.4u
m8815 4475 4388 71959 VSS nch l=0.04u w=0.8u
m8816 4476 4388 71960 VSS nch l=0.04u w=0.8u
m8817 4477 4388 71961 VSS nch l=0.04u w=0.8u
m8818 4478 4388 71962 VSS nch l=0.04u w=0.8u
m8819 4479 4388 71963 VSS nch l=0.04u w=0.8u
m8820 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8821 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8822 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8823 71964 4502 VSS VSS nch l=0.04u w=0.8u
m8824 71965 4503 VSS VSS nch l=0.04u w=0.8u
m8825 71966 4469 VSS VSS nch l=0.04u w=0.8u
m8826 71967 4470 VSS VSS nch l=0.04u w=0.8u
m8827 71968 4471 VSS VSS nch l=0.04u w=0.8u
m8828 71969 4472 VSS VSS nch l=0.04u w=0.8u
m8829 71970 4473 VSS VSS nch l=0.04u w=0.8u
m8830 4480 2427 71964 VSS nch l=0.04u w=0.8u
m8831 4481 4401 71965 VSS nch l=0.04u w=0.8u
m8832 4482 4458 71966 VSS nch l=0.04u w=0.8u
m8833 4483 4459 71967 VSS nch l=0.04u w=0.8u
m8834 4484 4460 71968 VSS nch l=0.04u w=0.8u
m8835 4485 4461 71969 VSS nch l=0.04u w=0.8u
m8836 4486 4462 71970 VSS nch l=0.04u w=0.8u
m8837 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8838 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8839 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8840 71971 2427 4480 VSS nch l=0.04u w=0.8u
m8841 71972 4401 4481 VSS nch l=0.04u w=0.8u
m8842 VSS 4502 71971 VSS nch l=0.04u w=0.8u
m8843 VSS 4503 71972 VSS nch l=0.04u w=0.8u
m8844 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8845 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8846 71973 4482 VSS VSS nch l=0.04u w=0.8u
m8847 71974 4483 VSS VSS nch l=0.04u w=0.8u
m8848 71975 4484 VSS VSS nch l=0.04u w=0.8u
m8849 71976 4485 VSS VSS nch l=0.04u w=0.8u
m8850 71977 4486 VSS VSS nch l=0.04u w=0.8u
m8851 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8852 4487 4475 71973 VSS nch l=0.04u w=0.8u
m8853 4488 4476 71974 VSS nch l=0.04u w=0.8u
m8854 4489 4477 71975 VSS nch l=0.04u w=0.8u
m8855 4490 4478 71976 VSS nch l=0.04u w=0.8u
m8856 4491 4479 71977 VSS nch l=0.04u w=0.8u
m8857 4493 2427 VSS VSS nch l=0.04u w=0.4u
m8858 4494 4401 VSS VSS nch l=0.04u w=0.4u
m8859 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8860 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8861 VSS 4452 VSS VSS nch l=0.26u w=0.8u
m8862 4496 4495 VSS VSS nch l=0.04u w=0.8u
m8863 4497 4487 VSS VSS nch l=0.04u w=0.4u
m8864 4498 4488 VSS VSS nch l=0.04u w=0.4u
m8865 4499 4489 VSS VSS nch l=0.04u w=0.4u
m8866 4500 4490 VSS VSS nch l=0.04u w=0.4u
m8867 4501 4491 VSS VSS nch l=0.04u w=0.4u
m8868 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8869 71978 4480 VSS VSS nch l=0.04u w=0.8u
m8870 71979 4481 VSS VSS nch l=0.04u w=0.8u
m8871 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8872 4502 4493 71978 VSS nch l=0.04u w=0.8u
m8873 4503 4494 71979 VSS nch l=0.04u w=0.8u
m8874 VSS 4505 4505 VSS nch l=0.04u w=0.8u
m8875 4506 4522 VSS VSS nch l=0.04u w=0.4u
m8876 4507 4523 VSS VSS nch l=0.04u w=0.4u
m8877 4508 4524 VSS VSS nch l=0.04u w=0.4u
m8878 4509 4525 VSS VSS nch l=0.04u w=0.4u
m8879 4510 4526 VSS VSS nch l=0.04u w=0.4u
m8880 VSS 4464 VSS VSS nch l=0.26u w=0.8u
m8881 VSS 4465 VSS VSS nch l=0.26u w=0.8u
m8882 71980 4493 4502 VSS nch l=0.04u w=0.8u
m8883 71981 4494 4503 VSS nch l=0.04u w=0.8u
m8884 VSS 4522 4506 VSS nch l=0.04u w=0.4u
m8885 VSS 4523 4507 VSS nch l=0.04u w=0.4u
m8886 VSS 4524 4508 VSS nch l=0.04u w=0.4u
m8887 VSS 4525 4509 VSS nch l=0.04u w=0.4u
m8888 VSS 4526 4510 VSS nch l=0.04u w=0.4u
m8889 4511 4512 VSS VSS nch l=0.04u w=0.8u
m8890 4514 4513 VSS VSS nch l=0.04u w=0.8u
m8891 VSS 4480 71980 VSS nch l=0.04u w=0.8u
m8892 VSS 4481 71981 VSS nch l=0.04u w=0.8u
m8893 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8894 4506 4522 VSS VSS nch l=0.04u w=0.4u
m8895 4507 4523 VSS VSS nch l=0.04u w=0.4u
m8896 4508 4524 VSS VSS nch l=0.04u w=0.4u
m8897 4509 4525 VSS VSS nch l=0.04u w=0.4u
m8898 4510 4526 VSS VSS nch l=0.04u w=0.4u
m8899 VSS 4522 4506 VSS nch l=0.04u w=0.4u
m8900 VSS 4523 4507 VSS nch l=0.04u w=0.4u
m8901 VSS 4524 4508 VSS nch l=0.04u w=0.4u
m8902 VSS 4525 4509 VSS nch l=0.04u w=0.4u
m8903 VSS 4526 4510 VSS nch l=0.04u w=0.4u
m8904 VSS 4515 4515 VSS nch l=0.04u w=0.8u
m8905 VSS 4518 4518 VSS nch l=0.04u w=0.8u
m8906 4520 4502 VSS VSS nch l=0.04u w=0.4u
m8907 4521 4503 VSS VSS nch l=0.04u w=0.4u
m8908 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8909 VSS 4502 4520 VSS nch l=0.04u w=0.4u
m8910 VSS 4503 4521 VSS nch l=0.04u w=0.4u
m8911 VSS 4527 4522 VSS nch l=0.04u w=0.4u
m8912 VSS 4528 4523 VSS nch l=0.04u w=0.4u
m8913 VSS 4529 4524 VSS nch l=0.04u w=0.4u
m8914 VSS 4530 4525 VSS nch l=0.04u w=0.4u
m8915 VSS 4531 4526 VSS nch l=0.04u w=0.4u
m8916 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m8917 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m8918 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8919 4520 4502 VSS VSS nch l=0.04u w=0.4u
m8920 4521 4503 VSS VSS nch l=0.04u w=0.4u
m8921 VSS 4502 4520 VSS nch l=0.04u w=0.4u
m8922 VSS 4503 4521 VSS nch l=0.04u w=0.4u
m8923 71982 4497 4527 VSS nch l=0.04u w=0.8u
m8924 71983 4498 4528 VSS nch l=0.04u w=0.8u
m8925 71984 4499 4529 VSS nch l=0.04u w=0.8u
m8926 71985 4500 4530 VSS nch l=0.04u w=0.8u
m8927 71986 4501 4531 VSS nch l=0.04u w=0.8u
m8928 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m8929 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m8930 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8931 VSS 4540 71982 VSS nch l=0.04u w=0.8u
m8932 VSS 4541 71983 VSS nch l=0.04u w=0.8u
m8933 VSS 4542 71984 VSS nch l=0.04u w=0.8u
m8934 VSS 4543 71985 VSS nch l=0.04u w=0.8u
m8935 VSS 4544 71986 VSS nch l=0.04u w=0.8u
m8936 4532 4520 VSS VSS nch l=0.04u w=0.4u
m8937 4533 4521 VSS VSS nch l=0.04u w=0.4u
m8938 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m8939 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m8940 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8941 VSS 4520 4532 VSS nch l=0.04u w=0.4u
m8942 VSS 4521 4533 VSS nch l=0.04u w=0.4u
m8943 4534 4497 VSS VSS nch l=0.04u w=0.4u
m8944 4535 4498 VSS VSS nch l=0.04u w=0.4u
m8945 4536 4499 VSS VSS nch l=0.04u w=0.4u
m8946 4537 4500 VSS VSS nch l=0.04u w=0.4u
m8947 4538 4501 VSS VSS nch l=0.04u w=0.4u
m8948 4532 4520 VSS VSS nch l=0.04u w=0.4u
m8949 4533 4521 VSS VSS nch l=0.04u w=0.4u
m8950 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m8951 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m8952 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8953 VSS 4520 4532 VSS nch l=0.04u w=0.4u
m8954 VSS 4521 4533 VSS nch l=0.04u w=0.4u
m8955 71987 4527 VSS VSS nch l=0.04u w=0.8u
m8956 71988 4528 VSS VSS nch l=0.04u w=0.8u
m8957 71989 4529 VSS VSS nch l=0.04u w=0.8u
m8958 71990 4530 VSS VSS nch l=0.04u w=0.8u
m8959 71991 4531 VSS VSS nch l=0.04u w=0.8u
m8960 4532 4520 VSS VSS nch l=0.04u w=0.4u
m8961 4533 4521 VSS VSS nch l=0.04u w=0.4u
m8962 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m8963 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m8964 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8965 4540 4534 71987 VSS nch l=0.04u w=0.8u
m8966 4541 4535 71988 VSS nch l=0.04u w=0.8u
m8967 4542 4536 71989 VSS nch l=0.04u w=0.8u
m8968 4543 4537 71990 VSS nch l=0.04u w=0.8u
m8969 4544 4538 71991 VSS nch l=0.04u w=0.8u
m8970 VSS 4520 4532 VSS nch l=0.04u w=0.4u
m8971 VSS 4521 4533 VSS nch l=0.04u w=0.4u
m8972 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m8973 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m8974 VSS 4504 VSS VSS nch l=0.26u w=0.8u
m8975 4545 4540 VSS VSS nch l=0.04u w=0.4u
m8976 4546 4541 VSS VSS nch l=0.04u w=0.4u
m8977 4547 4542 VSS VSS nch l=0.04u w=0.4u
m8978 4548 4543 VSS VSS nch l=0.04u w=0.4u
m8979 4549 4544 VSS VSS nch l=0.04u w=0.4u
m8980 4532 4520 VSS VSS nch l=0.04u w=0.4u
m8981 4533 4521 VSS VSS nch l=0.04u w=0.4u
m8982 4551 4550 VSS VSS nch l=0.04u w=0.8u
m8983 VSS 4520 4532 VSS nch l=0.04u w=0.4u
m8984 VSS 4521 4533 VSS nch l=0.04u w=0.4u
m8985 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m8986 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m8987 4554 4545 VSS VSS nch l=0.04u w=0.4u
m8988 4555 4546 VSS VSS nch l=0.04u w=0.4u
m8989 4556 4547 VSS VSS nch l=0.04u w=0.4u
m8990 4557 4548 VSS VSS nch l=0.04u w=0.4u
m8991 4558 4549 VSS VSS nch l=0.04u w=0.4u
m8992 4532 4520 VSS VSS nch l=0.04u w=0.4u
m8993 4533 4521 VSS VSS nch l=0.04u w=0.4u
m8994 VSS 4553 4553 VSS nch l=0.04u w=0.8u
m8995 VSS 4545 4554 VSS nch l=0.04u w=0.4u
m8996 VSS 4546 4555 VSS nch l=0.04u w=0.4u
m8997 VSS 4547 4556 VSS nch l=0.04u w=0.4u
m8998 VSS 4548 4557 VSS nch l=0.04u w=0.4u
m8999 VSS 4549 4558 VSS nch l=0.04u w=0.4u
m9000 VSS 4520 4532 VSS nch l=0.04u w=0.4u
m9001 VSS 4521 4533 VSS nch l=0.04u w=0.4u
m9002 VSS 4516 VSS VSS nch l=0.26u w=0.8u
m9003 VSS 4517 VSS VSS nch l=0.26u w=0.8u
m9004 4554 4545 VSS VSS nch l=0.04u w=0.4u
m9005 4555 4546 VSS VSS nch l=0.04u w=0.4u
m9006 4556 4547 VSS VSS nch l=0.04u w=0.4u
m9007 4557 4548 VSS VSS nch l=0.04u w=0.4u
m9008 4558 4549 VSS VSS nch l=0.04u w=0.4u
m9009 4532 4520 VSS VSS nch l=0.04u w=0.4u
m9010 4533 4521 VSS VSS nch l=0.04u w=0.4u
m9011 4559 4560 VSS VSS nch l=0.04u w=0.8u
m9012 4562 4561 VSS VSS nch l=0.04u w=0.8u
m9013 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9014 VSS 4545 4554 VSS nch l=0.04u w=0.4u
m9015 VSS 4546 4555 VSS nch l=0.04u w=0.4u
m9016 VSS 4547 4556 VSS nch l=0.04u w=0.4u
m9017 VSS 4548 4557 VSS nch l=0.04u w=0.4u
m9018 VSS 4549 4558 VSS nch l=0.04u w=0.4u
m9019 VSS 4520 4532 VSS nch l=0.04u w=0.4u
m9020 VSS 4521 4533 VSS nch l=0.04u w=0.4u
m9021 VSS 4564 4564 VSS nch l=0.04u w=0.8u
m9022 VSS 4567 4567 VSS nch l=0.04u w=0.8u
m9023 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9024 71992 4395 VSS VSS nch l=0.04u w=0.8u
m9025 71993 4395 VSS VSS nch l=0.04u w=0.8u
m9026 71994 4395 VSS VSS nch l=0.04u w=0.8u
m9027 71995 4395 VSS VSS nch l=0.04u w=0.8u
m9028 71996 4395 VSS VSS nch l=0.04u w=0.8u
m9029 4573 4606 VSS VSS nch l=0.04u w=0.4u
m9030 4574 4607 VSS VSS nch l=0.04u w=0.4u
m9031 4568 2666 71992 VSS nch l=0.04u w=0.8u
m9032 4569 2927 71993 VSS nch l=0.04u w=0.8u
m9033 4570 3205 71994 VSS nch l=0.04u w=0.8u
m9034 4571 4425 71995 VSS nch l=0.04u w=0.8u
m9035 4572 3937 71996 VSS nch l=0.04u w=0.8u
m9036 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9037 VSS 4606 4573 VSS nch l=0.04u w=0.4u
m9038 VSS 4607 4574 VSS nch l=0.04u w=0.4u
m9039 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9040 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9041 4573 4606 VSS VSS nch l=0.04u w=0.4u
m9042 4574 4607 VSS VSS nch l=0.04u w=0.4u
m9043 4575 DACPD VSS VSS nch l=0.04u w=0.4u
m9044 4576 DACPD VSS VSS nch l=0.04u w=0.4u
m9045 4577 DACPD VSS VSS nch l=0.04u w=0.4u
m9046 4578 DACPD VSS VSS nch l=0.04u w=0.4u
m9047 4579 DACPD VSS VSS nch l=0.04u w=0.4u
m9048 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9049 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9050 VSS 4606 4573 VSS nch l=0.04u w=0.4u
m9051 VSS 4607 4574 VSS nch l=0.04u w=0.4u
m9052 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9053 4573 4606 VSS VSS nch l=0.04u w=0.4u
m9054 4574 4607 VSS VSS nch l=0.04u w=0.4u
m9055 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9056 71997 DACPD VSS VSS nch l=0.04u w=0.8u
m9057 71998 DACPD VSS VSS nch l=0.04u w=0.8u
m9058 71999 DACPD VSS VSS nch l=0.04u w=0.8u
m9059 72000 DACPD VSS VSS nch l=0.04u w=0.8u
m9060 72001 DACPD VSS VSS nch l=0.04u w=0.8u
m9061 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9062 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9063 VSS 4606 4573 VSS nch l=0.04u w=0.4u
m9064 VSS 4607 4574 VSS nch l=0.04u w=0.4u
m9065 4580 DACPD 71997 VSS nch l=0.04u w=0.8u
m9066 4581 DACPD 71998 VSS nch l=0.04u w=0.8u
m9067 4582 DACPD 71999 VSS nch l=0.04u w=0.8u
m9068 4583 DACPD 72000 VSS nch l=0.04u w=0.8u
m9069 4584 DACPD 72001 VSS nch l=0.04u w=0.8u
m9070 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9071 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9072 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9073 4573 4606 VSS VSS nch l=0.04u w=0.4u
m9074 4574 4607 VSS VSS nch l=0.04u w=0.4u
m9075 72002 4575 VSS VSS nch l=0.04u w=0.8u
m9076 72003 4576 VSS VSS nch l=0.04u w=0.8u
m9077 72004 4577 VSS VSS nch l=0.04u w=0.8u
m9078 72005 4578 VSS VSS nch l=0.04u w=0.8u
m9079 72006 4579 VSS VSS nch l=0.04u w=0.8u
m9080 VSS 4606 4573 VSS nch l=0.04u w=0.4u
m9081 VSS 4607 4574 VSS nch l=0.04u w=0.4u
m9082 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9083 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9084 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9085 4586 4568 72002 VSS nch l=0.04u w=0.8u
m9086 4587 4569 72003 VSS nch l=0.04u w=0.8u
m9087 4588 4570 72004 VSS nch l=0.04u w=0.8u
m9088 4589 4571 72005 VSS nch l=0.04u w=0.8u
m9089 4590 4572 72006 VSS nch l=0.04u w=0.8u
m9090 4573 4606 VSS VSS nch l=0.04u w=0.4u
m9091 4574 4607 VSS VSS nch l=0.04u w=0.4u
m9092 VSS 4606 4573 VSS nch l=0.04u w=0.4u
m9093 VSS 4607 4574 VSS nch l=0.04u w=0.4u
m9094 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9095 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9096 VSS 4552 VSS VSS nch l=0.26u w=0.8u
m9097 72007 4586 VSS VSS nch l=0.04u w=0.8u
m9098 72008 4587 VSS VSS nch l=0.04u w=0.8u
m9099 72009 4588 VSS VSS nch l=0.04u w=0.8u
m9100 72010 4589 VSS VSS nch l=0.04u w=0.8u
m9101 72011 4590 VSS VSS nch l=0.04u w=0.8u
m9102 4573 4606 VSS VSS nch l=0.04u w=0.4u
m9103 4574 4607 VSS VSS nch l=0.04u w=0.4u
m9104 4597 4596 VSS VSS nch l=0.04u w=0.8u
m9105 4591 4580 72007 VSS nch l=0.04u w=0.8u
m9106 4592 4581 72008 VSS nch l=0.04u w=0.8u
m9107 4593 4582 72009 VSS nch l=0.04u w=0.8u
m9108 4594 4583 72010 VSS nch l=0.04u w=0.8u
m9109 4595 4584 72011 VSS nch l=0.04u w=0.8u
m9110 VSS 4606 4573 VSS nch l=0.04u w=0.4u
m9111 VSS 4607 4574 VSS nch l=0.04u w=0.4u
m9112 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9113 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9114 VSS 4599 4599 VSS nch l=0.04u w=0.8u
m9115 4601 155 VSS VSS nch l=0.04u w=0.4u
m9116 4602 155 VSS VSS nch l=0.04u w=0.4u
m9117 4603 155 VSS VSS nch l=0.04u w=0.4u
m9118 4604 155 VSS VSS nch l=0.04u w=0.4u
m9119 4605 155 VSS VSS nch l=0.04u w=0.4u
m9120 4606 4624 VSS VSS nch l=0.04u w=0.4u
m9121 4607 4625 VSS VSS nch l=0.04u w=0.4u
m9122 VSS 4565 VSS VSS nch l=0.26u w=0.8u
m9123 VSS 4566 VSS VSS nch l=0.26u w=0.8u
m9124 VSS 4624 4606 VSS nch l=0.04u w=0.4u
m9125 VSS 4625 4607 VSS nch l=0.04u w=0.4u
m9126 4608 4609 VSS VSS nch l=0.04u w=0.8u
m9127 4611 4610 VSS VSS nch l=0.04u w=0.8u
m9128 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9129 72012 155 VSS VSS nch l=0.04u w=0.8u
m9130 72013 155 VSS VSS nch l=0.04u w=0.8u
m9131 72014 155 VSS VSS nch l=0.04u w=0.8u
m9132 72015 155 VSS VSS nch l=0.04u w=0.8u
m9133 72016 155 VSS VSS nch l=0.04u w=0.8u
m9134 4606 4624 VSS VSS nch l=0.04u w=0.4u
m9135 4607 4625 VSS VSS nch l=0.04u w=0.4u
m9136 4612 4392 72012 VSS nch l=0.04u w=0.8u
m9137 4613 4392 72013 VSS nch l=0.04u w=0.8u
m9138 4614 4392 72014 VSS nch l=0.04u w=0.8u
m9139 4615 4392 72015 VSS nch l=0.04u w=0.8u
m9140 4616 4392 72016 VSS nch l=0.04u w=0.8u
m9141 VSS 4624 4606 VSS nch l=0.04u w=0.4u
m9142 VSS 4625 4607 VSS nch l=0.04u w=0.4u
m9143 4617 4649 VSS VSS nch l=0.04u w=0.4u
m9144 FOUTVCO 4639 VSS VSS nch l=0.04u w=0.4u
m9145 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9146 VSS 4649 4617 VSS nch l=0.04u w=0.4u
m9147 VSS 4639 FOUTVCO VSS nch l=0.04u w=0.4u
m9148 72017 4601 VSS VSS nch l=0.04u w=0.8u
m9149 72018 4602 VSS VSS nch l=0.04u w=0.8u
m9150 72019 4603 VSS VSS nch l=0.04u w=0.8u
m9151 72020 4604 VSS VSS nch l=0.04u w=0.8u
m9152 72021 4605 VSS VSS nch l=0.04u w=0.8u
m9153 72022 4640 VSS VSS nch l=0.04u w=0.8u
m9154 72023 4641 VSS VSS nch l=0.04u w=0.8u
m9155 4617 4649 VSS VSS nch l=0.04u w=0.4u
m9156 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9157 FOUTVCO 4639 VSS VSS nch l=0.04u w=0.4u
m9158 4619 4591 72017 VSS nch l=0.04u w=0.8u
m9159 4620 4592 72018 VSS nch l=0.04u w=0.8u
m9160 4621 4593 72019 VSS nch l=0.04u w=0.8u
m9161 4622 4594 72020 VSS nch l=0.04u w=0.8u
m9162 4623 4595 72021 VSS nch l=0.04u w=0.8u
m9163 4624 2426 72022 VSS nch l=0.04u w=0.8u
m9164 4625 4426 72023 VSS nch l=0.04u w=0.8u
m9165 VSS 4649 4617 VSS nch l=0.04u w=0.4u
m9166 VSS 4639 FOUTVCO VSS nch l=0.04u w=0.4u
m9167 72024 2426 4624 VSS nch l=0.04u w=0.8u
m9168 72025 4426 4625 VSS nch l=0.04u w=0.8u
m9169 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9170 4617 4649 VSS VSS nch l=0.04u w=0.4u
m9171 FOUTVCO 4639 VSS VSS nch l=0.04u w=0.4u
m9172 VSS 4640 72024 VSS nch l=0.04u w=0.8u
m9173 VSS 4641 72025 VSS nch l=0.04u w=0.8u
m9174 72026 4619 VSS VSS nch l=0.04u w=0.8u
m9175 72027 4620 VSS VSS nch l=0.04u w=0.8u
m9176 72028 4621 VSS VSS nch l=0.04u w=0.8u
m9177 72029 4622 VSS VSS nch l=0.04u w=0.8u
m9178 72030 4623 VSS VSS nch l=0.04u w=0.8u
m9179 VSS 4649 4617 VSS nch l=0.04u w=0.4u
m9180 VSS 4639 FOUTVCO VSS nch l=0.04u w=0.4u
m9181 4627 4612 72026 VSS nch l=0.04u w=0.8u
m9182 4628 4613 72027 VSS nch l=0.04u w=0.8u
m9183 4629 4614 72028 VSS nch l=0.04u w=0.8u
m9184 4630 4615 72029 VSS nch l=0.04u w=0.8u
m9185 4631 4616 72030 VSS nch l=0.04u w=0.8u
m9186 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9187 4617 4649 VSS VSS nch l=0.04u w=0.4u
m9188 FOUTVCO 4639 VSS VSS nch l=0.04u w=0.4u
m9189 4632 2426 VSS VSS nch l=0.04u w=0.4u
m9190 4633 4426 VSS VSS nch l=0.04u w=0.4u
m9191 VSS 4649 4617 VSS nch l=0.04u w=0.4u
m9192 VSS 4639 FOUTVCO VSS nch l=0.04u w=0.4u
m9193 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9194 4634 4627 VSS VSS nch l=0.04u w=0.4u
m9195 4635 4628 VSS VSS nch l=0.04u w=0.4u
m9196 4636 4629 VSS VSS nch l=0.04u w=0.4u
m9197 4637 4630 VSS VSS nch l=0.04u w=0.4u
m9198 4638 4631 VSS VSS nch l=0.04u w=0.4u
m9199 72031 4624 VSS VSS nch l=0.04u w=0.8u
m9200 72032 4625 VSS VSS nch l=0.04u w=0.8u
m9201 4642 4649 VSS VSS nch l=0.04u w=0.4u
m9202 4643 4642 4639 VSS nch l=0.04u w=0.8u
m9203 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9204 4640 4632 72031 VSS nch l=0.04u w=0.8u
m9205 4641 4633 72032 VSS nch l=0.04u w=0.8u
m9206 4644 4659 VSS VSS nch l=0.04u w=0.4u
m9207 4645 4660 VSS VSS nch l=0.04u w=0.4u
m9208 4646 4661 VSS VSS nch l=0.04u w=0.4u
m9209 4647 4662 VSS VSS nch l=0.04u w=0.4u
m9210 4648 4663 VSS VSS nch l=0.04u w=0.4u
m9211 VSS 4649 4642 VSS nch l=0.04u w=0.4u
m9212 VSS 4687 4643 VSS nch l=0.04u w=0.8u
m9213 72033 4632 4640 VSS nch l=0.04u w=0.8u
m9214 72034 4633 4641 VSS nch l=0.04u w=0.8u
m9215 VSS 4659 4644 VSS nch l=0.04u w=0.4u
m9216 VSS 4660 4645 VSS nch l=0.04u w=0.4u
m9217 VSS 4661 4646 VSS nch l=0.04u w=0.4u
m9218 VSS 4662 4647 VSS nch l=0.04u w=0.4u
m9219 VSS 4663 4648 VSS nch l=0.04u w=0.4u
m9220 4643 4687 VSS VSS nch l=0.04u w=0.8u
m9221 VSS 4598 VSS VSS nch l=0.26u w=0.8u
m9222 VSS 4624 72033 VSS nch l=0.04u w=0.8u
m9223 VSS 4625 72034 VSS nch l=0.04u w=0.8u
m9224 4644 4659 VSS VSS nch l=0.04u w=0.4u
m9225 4645 4660 VSS VSS nch l=0.04u w=0.4u
m9226 4646 4661 VSS VSS nch l=0.04u w=0.4u
m9227 4647 4662 VSS VSS nch l=0.04u w=0.4u
m9228 4648 4663 VSS VSS nch l=0.04u w=0.4u
m9229 4649 4679 VSS VSS nch l=0.04u w=0.4u
m9230 4652 4651 VSS VSS nch l=0.04u w=0.8u
m9231 VSS 4659 4644 VSS nch l=0.04u w=0.4u
m9232 VSS 4660 4645 VSS nch l=0.04u w=0.4u
m9233 VSS 4661 4646 VSS nch l=0.04u w=0.4u
m9234 VSS 4662 4647 VSS nch l=0.04u w=0.4u
m9235 VSS 4663 4648 VSS nch l=0.04u w=0.4u
m9236 VSS 4679 4649 VSS nch l=0.04u w=0.4u
m9237 VSS 4699 4650 VSS nch l=0.04u w=0.8u
m9238 4657 4640 VSS VSS nch l=0.04u w=0.4u
m9239 4658 4641 VSS VSS nch l=0.04u w=0.4u
m9240 4649 4679 VSS VSS nch l=0.04u w=0.4u
m9241 4650 4699 VSS VSS nch l=0.04u w=0.8u
m9242 VSS 4656 4656 VSS nch l=0.04u w=0.8u
m9243 VSS 4640 4657 VSS nch l=0.04u w=0.4u
m9244 VSS 4641 4658 VSS nch l=0.04u w=0.4u
m9245 VSS 4664 4659 VSS nch l=0.04u w=0.4u
m9246 VSS 4665 4660 VSS nch l=0.04u w=0.4u
m9247 VSS 4666 4661 VSS nch l=0.04u w=0.4u
m9248 VSS 4667 4662 VSS nch l=0.04u w=0.4u
m9249 VSS 4668 4663 VSS nch l=0.04u w=0.4u
m9250 VSS 4679 4649 VSS nch l=0.04u w=0.4u
m9251 4654 4642 4650 VSS nch l=0.04u w=0.8u
m9252 4657 4640 VSS VSS nch l=0.04u w=0.4u
m9253 4658 4641 VSS VSS nch l=0.04u w=0.4u
m9254 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9255 VSS 4640 4657 VSS nch l=0.04u w=0.4u
m9256 VSS 4641 4658 VSS nch l=0.04u w=0.4u
m9257 72035 4634 4664 VSS nch l=0.04u w=0.8u
m9258 72036 4635 4665 VSS nch l=0.04u w=0.8u
m9259 72037 4636 4666 VSS nch l=0.04u w=0.8u
m9260 72038 4637 4667 VSS nch l=0.04u w=0.8u
m9261 72039 4638 4668 VSS nch l=0.04u w=0.8u
m9262 4669 4654 VSS VSS nch l=0.04u w=0.4u
m9263 VSS 4682 72035 VSS nch l=0.04u w=0.8u
m9264 VSS 4683 72036 VSS nch l=0.04u w=0.8u
m9265 VSS 4684 72037 VSS nch l=0.04u w=0.8u
m9266 VSS 4685 72038 VSS nch l=0.04u w=0.8u
m9267 VSS 4686 72039 VSS nch l=0.04u w=0.8u
m9268 VSS 4654 4669 VSS nch l=0.04u w=0.4u
m9269 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9270 4671 4657 VSS VSS nch l=0.04u w=0.4u
m9271 4672 4658 VSS VSS nch l=0.04u w=0.4u
m9272 VSS PD 4670 VSS nch l=0.04u w=0.15u
m9273 4669 4654 VSS VSS nch l=0.04u w=0.4u
m9274 VSS 4657 4671 VSS nch l=0.04u w=0.4u
m9275 VSS 4658 4672 VSS nch l=0.04u w=0.4u
m9276 4673 PD VSS VSS nch l=0.04u w=0.15u
m9277 4674 4634 VSS VSS nch l=0.04u w=0.4u
m9278 4675 4635 VSS VSS nch l=0.04u w=0.4u
m9279 4676 4636 VSS VSS nch l=0.04u w=0.4u
m9280 4677 4637 VSS VSS nch l=0.04u w=0.4u
m9281 4678 4638 VSS VSS nch l=0.04u w=0.4u
m9282 VSS 4654 4669 VSS nch l=0.04u w=0.4u
m9283 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9284 4671 4657 VSS VSS nch l=0.04u w=0.4u
m9285 4672 4658 VSS VSS nch l=0.04u w=0.4u
m9286 4669 4654 VSS VSS nch l=0.04u w=0.4u
m9287 VSS 4657 4671 VSS nch l=0.04u w=0.4u
m9288 VSS 4658 4672 VSS nch l=0.04u w=0.4u
m9289 VSS 4654 4669 VSS nch l=0.04u w=0.4u
m9290 72041 4664 VSS VSS nch l=0.04u w=0.8u
m9291 72042 4665 VSS VSS nch l=0.04u w=0.8u
m9292 72043 4666 VSS VSS nch l=0.04u w=0.8u
m9293 72044 4667 VSS VSS nch l=0.04u w=0.8u
m9294 72045 4668 VSS VSS nch l=0.04u w=0.8u
m9295 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9296 VSS 4680 4680 VSS nch l=0.04u w=0.8u
m9297 4671 4657 VSS VSS nch l=0.04u w=0.4u
m9298 4672 4658 VSS VSS nch l=0.04u w=0.4u
m9299 4669 4654 VSS VSS nch l=0.04u w=0.4u
m9300 4682 4674 72041 VSS nch l=0.04u w=0.8u
m9301 4683 4675 72042 VSS nch l=0.04u w=0.8u
m9302 4684 4676 72043 VSS nch l=0.04u w=0.8u
m9303 4685 4677 72044 VSS nch l=0.04u w=0.8u
m9304 4686 4678 72045 VSS nch l=0.04u w=0.8u
m9305 4679 4673 VSS VSS nch l=0.04u w=0.8u
m9306 VSS 4657 4671 VSS nch l=0.04u w=0.4u
m9307 VSS 4658 4672 VSS nch l=0.04u w=0.4u
m9308 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9309 VSS 4654 4669 VSS nch l=0.04u w=0.4u
m9310 VSS 4673 4679 VSS nch l=0.04u w=0.8u
m9311 4688 4682 VSS VSS nch l=0.04u w=0.4u
m9312 4689 4683 VSS VSS nch l=0.04u w=0.4u
m9313 4690 4684 VSS VSS nch l=0.04u w=0.4u
m9314 4691 4685 VSS VSS nch l=0.04u w=0.4u
m9315 4692 4686 VSS VSS nch l=0.04u w=0.4u
m9316 4671 4657 VSS VSS nch l=0.04u w=0.4u
m9317 4672 4658 VSS VSS nch l=0.04u w=0.4u
m9318 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9319 4687 FOUTVCOPD VSS VSS nch l=0.04u w=0.4u
m9320 VSS 4670 4693 VSS nch l=0.04u w=0.8u
m9321 VSS 4657 4671 VSS nch l=0.04u w=0.4u
m9322 VSS 4658 4672 VSS nch l=0.04u w=0.4u
m9323 VSS PD 4687 VSS nch l=0.04u w=0.4u
m9324 4694 4688 VSS VSS nch l=0.04u w=0.4u
m9325 4695 4689 VSS VSS nch l=0.04u w=0.4u
m9326 4696 4690 VSS VSS nch l=0.04u w=0.4u
m9327 4697 4691 VSS VSS nch l=0.04u w=0.4u
m9328 4698 4692 VSS VSS nch l=0.04u w=0.4u
m9329 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9330 4671 4657 VSS VSS nch l=0.04u w=0.4u
m9331 4672 4658 VSS VSS nch l=0.04u w=0.4u
m9332 VSS 4688 4694 VSS nch l=0.04u w=0.4u
m9333 VSS 4689 4695 VSS nch l=0.04u w=0.4u
m9334 VSS 4690 4696 VSS nch l=0.04u w=0.4u
m9335 VSS 4691 4697 VSS nch l=0.04u w=0.4u
m9336 VSS 4692 4698 VSS nch l=0.04u w=0.4u
m9337 VSS 4657 4671 VSS nch l=0.04u w=0.4u
m9338 VSS 4658 4672 VSS nch l=0.04u w=0.4u
m9339 4699 PD VSS VSS nch l=0.04u w=0.4u
m9340 4694 4688 VSS VSS nch l=0.04u w=0.4u
m9341 4695 4689 VSS VSS nch l=0.04u w=0.4u
m9342 4696 4690 VSS VSS nch l=0.04u w=0.4u
m9343 4697 4691 VSS VSS nch l=0.04u w=0.4u
m9344 4698 4692 VSS VSS nch l=0.04u w=0.4u
m9345 VSS 4655 VSS VSS nch l=0.26u w=0.8u
m9346 4671 4657 VSS VSS nch l=0.04u w=0.4u
m9347 4672 4658 VSS VSS nch l=0.04u w=0.4u
m9348 VSS FOUTPOSTDIVPD 4699 VSS nch l=0.04u w=0.4u
m9349 VSS 4688 4694 VSS nch l=0.04u w=0.4u
m9350 VSS 4689 4695 VSS nch l=0.04u w=0.4u
m9351 VSS 4690 4696 VSS nch l=0.04u w=0.4u
m9352 VSS 4691 4697 VSS nch l=0.04u w=0.4u
m9353 VSS 4692 4698 VSS nch l=0.04u w=0.4u
m9354 4702 4701 VSS VSS nch l=0.04u w=0.8u
m9355 VSS 4657 4671 VSS nch l=0.04u w=0.4u
m9356 VSS 4658 4672 VSS nch l=0.04u w=0.4u
m9357 4703 FOUTPOSTDIVPD VSS VSS nch l=0.04u w=0.4u
m9358 72081 4703 VSS VSS nch l=0.04u w=0.8u
m9359 4705 4669 VSS VSS nch l=0.04u w=0.4u
m9360 4704 12 72081 VSS nch l=0.04u w=0.8u
m9361 VSS 4669 4705 VSS nch l=0.04u w=0.4u
m9362 4673 4670 VSS VSS nch l=0.04u w=0.4u
m9363 4707 4704 VSS VSS nch l=0.04u w=0.4u
m9364 VSS 4788 4706 VSS nch l=0.04u w=0.8u
m9365 VSS 4670 4673 VSS nch l=0.04u w=0.4u
m9366 VSS 4704 4707 VSS nch l=0.04u w=0.4u
m9367 4706 4788 VSS VSS nch l=0.04u w=0.8u
m9368 VSS 4788 4706 VSS nch l=0.04u w=0.8u
m9369 4670 4929 VSS VSS nch l=0.04u w=0.4u
m9370 4706 4788 VSS VSS nch l=0.04u w=0.8u
m9371 4709 POSTDIV2[1] VSS VSS nch l=0.04u w=0.4u
m9372 VSS 4929 4670 VSS nch l=0.04u w=0.4u
m9373 VSS 4788 4706 VSS nch l=0.04u w=0.8u
m9374 VSS POSTDIV2[2] 4709 VSS nch l=0.04u w=0.4u
m9375 4706 4788 VSS VSS nch l=0.04u w=0.8u
m9376 VSS 4788 4706 VSS nch l=0.04u w=0.8u
m9377 4710 4709 VSS VSS nch l=0.04u w=0.4u
m9378 4706 4788 VSS VSS nch l=0.04u w=0.8u
m9379 4708 4669 4706 VSS nch l=0.04u w=0.8u
m9380 4711 4860 VSS VSS nch l=0.04u w=0.4u
m9381 VSS VSS VSS VSS nch l=0.19u w=2.6u
m9382 4706 4669 4708 VSS nch l=0.04u w=0.8u
m9383 VSS 4710 4711 VSS nch l=0.04u w=0.4u
m9384 72115 4929 VSS VSS nch l=0.19u w=2.6u
m9385 4708 4669 4706 VSS nch l=0.04u w=0.8u
m9386 4713 4953 VSS VSS nch l=0.04u w=0.4u
m9387 72117 POSTDIV2[0] VSS VSS nch l=0.04u w=0.8u
m9388 4712 4929 72115 VSS nch l=0.19u w=2.6u
m9389 4715 POSTDIV1[1] VSS VSS nch l=0.04u w=0.4u
m9390 4714 POSTDIV2[1] 72117 VSS nch l=0.04u w=0.8u
m9391 72120 4929 4712 VSS nch l=0.19u w=2.6u
m9392 VSS POSTDIV1[2] 4715 VSS nch l=0.04u w=0.4u
m9393 VSS 4787 4716 VSS nch l=0.04u w=0.4u
m9394 4786 POSTDIV2[0] VSS VSS nch l=0.04u w=0.4u
m9395 VSS 4929 72120 VSS nch l=0.19u w=2.6u
m9396 72123 4709 VSS VSS nch l=0.04u w=0.8u
m9397 VSS POSTDIV2[1] 4786 VSS nch l=0.04u w=0.4u
m9398 72124 4790 4787 VSS nch l=0.04u w=0.8u
m9399 4788 4715 72123 VSS nch l=0.04u w=0.8u
m9400 72125 4929 VSS VSS nch l=0.19u w=2.6u
m9401 VSS 4713 72124 VSS nch l=0.04u w=0.8u
m9402 4789 POSTDIV2[2] VSS VSS nch l=0.04u w=0.4u
m9403 4712 4929 72125 VSS nch l=0.19u w=2.6u
m9404 4791 4860 VSS VSS nch l=0.04u w=0.4u
m9405 VSS 4793 4790 VSS nch l=0.04u w=0.4u
m9406 VSS 4788 4791 VSS nch l=0.04u w=0.4u
m9407 72129 4929 4712 VSS nch l=0.19u w=2.6u
m9408 4792 4789 VSS VSS nch l=0.04u w=0.4u
m9409 72130 4716 VSS VSS nch l=0.04u w=0.12u
m9410 VSS 4714 4792 VSS nch l=0.04u w=0.4u
m9411 VSS 4929 72129 VSS nch l=0.19u w=2.6u
m9412 4793 4874 72130 VSS nch l=0.04u w=0.12u
m9413 4794 BYPASS VSS VSS nch l=0.04u w=0.4u
m9414 4857 4981 4793 VSS nch l=0.04u w=0.4u
m9415 VSS FOUTPOSTDIVPD 4794 VSS nch l=0.04u w=0.4u
m9416 72135 4929 VSS VSS nch l=0.19u w=2.6u
m9417 72136 4789 VSS VSS nch l=0.04u w=0.8u
m9418 4858 4714 72136 VSS nch l=0.04u w=0.8u
m9419 4712 4929 72135 VSS nch l=0.19u w=2.6u
m9420 72138 4870 4857 VSS nch l=0.04u w=0.8u
m9421 4860 4794 VSS VSS nch l=0.04u w=0.4u
m9422 VSS 4713 72138 VSS nch l=0.04u w=0.8u
m9423 4863 4789 VSS VSS nch l=0.04u w=0.4u
m9424 72142 4929 4712 VSS nch l=0.19u w=2.6u
m9425 72143 4857 VSS VSS nch l=0.04u w=0.24u
m9426 4866 POSTDIV1[0] VSS VSS nch l=0.04u w=0.4u
m9427 VSS 4786 4863 VSS nch l=0.04u w=0.4u
m9428 4870 4981 72143 VSS nch l=0.04u w=0.24u
m9429 VSS 4929 72142 VSS nch l=0.19u w=2.6u
m9430 4871 4874 4870 VSS nch l=0.04u w=0.4u
m9431 4872 POSTDIV1[1] VSS VSS nch l=0.04u w=0.4u
m9432 4873 POSTDIV2[1] VSS VSS nch l=0.04u w=0.4u
m9433 72146 4929 VSS VSS nch l=0.19u w=2.6u
m9434 4874 4981 VSS VSS nch l=0.04u w=0.4u
m9435 4712 4929 72146 VSS nch l=0.19u w=2.6u
m9436 4875 POSTDIV1[2] VSS VSS nch l=0.04u w=0.4u
m9437 4876 POSTDIV2[0] VSS VSS nch l=0.04u w=0.4u
m9438 VSS 4873 4876 VSS nch l=0.04u w=0.4u
m9439 72150 4929 4712 VSS nch l=0.19u w=2.6u
m9440 VSS 4926 4871 VSS nch l=0.04u w=0.4u
m9441 4925 POSTDIV1[0] VSS VSS nch l=0.04u w=0.4u
m9442 4876 4789 VSS VSS nch l=0.04u w=0.4u
m9443 VSS 4929 72150 VSS nch l=0.19u w=2.6u
m9444 VSS 4872 4925 VSS nch l=0.04u w=0.4u
m9445 4925 POSTDIV1[2] VSS VSS nch l=0.04u w=0.4u
m9446 72154 4931 4926 VSS nch l=0.04u w=0.8u
m9447 VSS 4792 4927 VSS nch l=0.04u w=0.8u
m9448 72155 4974 VSS VSS nch l=0.19u w=2.6u
m9449 VSS 4713 72154 VSS nch l=0.04u w=0.8u
m9450 4927 4792 VSS VSS nch l=0.04u w=0.8u
m9451 4929 4974 72155 VSS nch l=0.19u w=2.6u
m9452 72157 4866 VSS VSS nch l=0.04u w=0.8u
m9453 4928 5527 4927 VSS nch l=0.04u w=0.8u
m9454 72159 4872 72157 VSS nch l=0.04u w=0.8u
m9455 VSS 4934 4931 VSS nch l=0.04u w=0.4u
m9456 72160 4974 4929 VSS nch l=0.19u w=2.6u
m9457 4930 POSTDIV1[2] 72159 VSS nch l=0.04u w=0.8u
m9458 72162 4871 VSS VSS nch l=0.04u w=0.12u
m9459 4932 4928 VSS VSS nch l=0.04u w=0.4u
m9460 4934 4951 72162 VSS nch l=0.04u w=0.12u
m9461 VSS 4974 72160 VSS nch l=0.19u w=2.6u
m9462 4936 4981 4934 VSS nch l=0.04u w=0.4u
m9463 72167 4930 4933 VSS nch l=0.04u w=0.8u
m9464 4937 4932 4935 VSS nch l=0.04u w=0.4u
m9465 72168 4974 VSS VSS nch l=0.19u w=2.6u
m9466 4938 4939 VSS VSS nch l=0.04u w=0.8u
m9467 VSS 4941 72167 VSS nch l=0.04u w=0.8u
m9468 72170 4928 4937 VSS nch l=0.04u w=0.12u
m9469 72171 4945 4936 VSS nch l=0.04u w=0.8u
m9470 4929 4974 72168 VSS nch l=0.19u w=2.6u
m9471 VSS 4942 72170 VSS nch l=0.04u w=0.12u
m9472 VSS PD 4940 VSS nch l=0.04u w=0.4u
m9473 VSS 4713 72171 VSS nch l=0.04u w=0.8u
m9474 72173 POSTDIV1[0] VSS VSS nch l=0.04u w=0.8u
m9475 4942 4937 VSS VSS nch l=0.04u w=0.4u
m9476 4943 4940 VSS VSS nch l=0.04u w=0.4u
m9477 72174 4974 4929 VSS nch l=0.19u w=2.6u
m9478 72175 4936 VSS VSS nch l=0.04u w=0.24u
m9479 72176 POSTDIV1[1] 72173 VSS nch l=0.04u w=0.8u
m9480 4944 FOUT4PHASEPD VSS VSS nch l=0.04u w=0.4u
m9481 4945 4981 72175 VSS nch l=0.04u w=0.24u
m9482 4941 4875 72176 VSS nch l=0.04u w=0.8u
m9483 VSS 4974 72174 VSS nch l=0.19u w=2.6u
m9484 4947 4928 4942 VSS nch l=0.04u w=0.4u
m9485 VSS FOUTPOSTDIVPD 4944 VSS nch l=0.04u w=0.4u
m9486 4713 4951 4945 VSS nch l=0.04u w=0.4u
m9487 72177 4932 4947 VSS nch l=0.04u w=0.12u
m9488 4944 PD VSS VSS nch l=0.04u w=0.4u
m9489 72179 4974 VSS VSS nch l=0.19u w=2.6u
m9490 72180 POSTDIV1[0] VSS VSS nch l=0.04u w=0.8u
m9491 VSS 4952 72177 VSS nch l=0.04u w=0.12u
m9492 4951 4981 VSS VSS nch l=0.04u w=0.4u
m9493 72183 4872 72180 VSS nch l=0.04u w=0.8u
m9494 4952 4947 VSS VSS nch l=0.04u w=0.4u
m9495 4929 4974 72179 VSS nch l=0.19u w=2.6u
m9496 4953 4944 VSS VSS nch l=0.04u w=0.4u
m9497 4950 POSTDIV1[2] 72183 VSS nch l=0.04u w=0.8u
m9498 72185 4974 4929 VSS nch l=0.19u w=2.6u
m9499 FOUT1PH270 4970 VSS VSS nch l=0.04u w=0.4u
m9500 4957 4958 VSS VSS nch l=0.04u w=0.8u
m9501 4959 4953 VSS VSS nch l=0.04u w=0.4u
m9502 4960 4792 VSS VSS nch l=0.04u w=0.4u
m9503 VSS 4970 FOUT1PH270 VSS nch l=0.04u w=0.4u
m9504 72186 4950 4956 VSS nch l=0.04u w=0.8u
m9505 VSS 4974 72185 VSS nch l=0.19u w=2.6u
m9506 FOUT1PH270 4970 VSS VSS nch l=0.04u w=0.4u
m9507 VSS 4968 72186 VSS nch l=0.04u w=0.8u
m9508 VSS 1580 4961 VSS nch l=0.04u w=0.4u
m9509 72188 4792 VSS VSS nch l=0.04u w=0.8u
m9510 VSS 4970 FOUT1PH270 VSS nch l=0.04u w=0.4u
m9511 72189 4974 VSS VSS nch l=0.19u w=2.6u
m9512 4964 4961 VSS VSS nch l=0.04u w=0.4u
m9513 VSS 4966 4962 VSS nch l=0.04u w=0.4u
m9514 4963 4952 72188 VSS nch l=0.04u w=0.8u
m9515 FOUT1PH270 4970 VSS VSS nch l=0.04u w=0.4u
m9516 4965 4968 VSS VSS nch l=0.04u w=0.4u
m9517 4929 4974 72189 VSS nch l=0.19u w=2.6u
m9518 VSS 4970 FOUT1PH270 VSS nch l=0.04u w=0.4u
m9519 72190 4969 4966 VSS nch l=0.04u w=0.8u
m9520 72191 4960 VSS VSS nch l=0.04u w=0.8u
m9521 FOUT1PH270 4970 VSS VSS nch l=0.04u w=0.4u
m9522 72192 4866 VSS VSS nch l=0.04u w=0.8u
m9523 72193 4974 4929 VSS nch l=0.19u w=2.6u
m9524 VSS 4959 72190 VSS nch l=0.04u w=0.8u
m9525 4967 4935 72191 VSS nch l=0.04u w=0.8u
m9526 VSS 4970 FOUT1PH270 VSS nch l=0.04u w=0.4u
m9527 72197 POSTDIV1[1] 72192 VSS nch l=0.04u w=0.8u
m9528 VSS 4974 72193 VSS nch l=0.19u w=2.6u
m9529 4968 POSTDIV1[2] 72197 VSS nch l=0.04u w=0.8u
m9530 VSS 4978 4969 VSS nch l=0.04u w=0.4u
m9531 72199 4967 VSS VSS nch l=0.04u w=0.8u
m9532 4973 5424 4970 VSS nch l=0.04u w=0.8u
m9533 72200 4712 VSS VSS nch l=0.19u w=2.6u
m9534 72201 4962 VSS VSS nch l=0.04u w=0.12u
m9535 4972 4963 72199 VSS nch l=0.04u w=0.8u
m9536 VSS 4716 4973 VSS nch l=0.04u w=0.8u
m9537 4975 4976 VSS VSS nch l=0.04u w=0.8u
m9538 4977 4866 VSS VSS nch l=0.04u w=0.4u
m9539 4978 4997 72201 VSS nch l=0.04u w=0.12u
m9540 4974 4712 72200 VSS nch l=0.19u w=2.6u
m9541 72202 4963 4972 VSS nch l=0.04u w=0.8u
m9542 4973 4716 VSS VSS nch l=0.04u w=0.8u
m9543 VSS 4872 4977 VSS nch l=0.04u w=0.4u
m9544 4980 5143 4978 VSS nch l=0.04u w=0.4u
m9545 VSS 4967 72202 VSS nch l=0.04u w=0.8u
m9546 VSS 1487 4979 VSS nch l=0.04u w=0.4u
m9547 4977 4875 VSS VSS nch l=0.04u w=0.4u
m9548 72203 4712 4974 VSS nch l=0.19u w=2.6u
m9549 VSS 4986 4981 VSS nch l=0.04u w=0.4u
m9550 4983 4979 VSS VSS nch l=0.04u w=0.4u
m9551 72204 4990 4980 VSS nch l=0.04u w=0.8u
m9552 VSS 4863 4982 VSS nch l=0.04u w=0.8u
m9553 4986 5424 VSS VSS nch l=0.04u w=0.4u
m9554 VSS 4712 72203 VSS nch l=0.19u w=2.6u
m9555 VSS 4977 4984 VSS nch l=0.04u w=0.8u
m9556 VSS 4959 72204 VSS nch l=0.04u w=0.8u
m9557 4982 4863 VSS VSS nch l=0.04u w=0.8u
m9558 4984 4977 VSS VSS nch l=0.04u w=0.8u
m9559 72205 4712 VSS VSS nch l=0.19u w=2.6u
m9560 72207 4980 VSS VSS nch l=0.04u w=0.24u
m9561 4985 5527 4982 VSS nch l=0.04u w=0.8u
m9562 4987 FOUT1PH270 VSS VSS nch l=0.04u w=0.4u
m9563 VSS 4977 4984 VSS nch l=0.04u w=0.8u
m9564 4990 5143 72207 VSS nch l=0.04u w=0.24u
m9565 VSS FOUT1PH270 4987 VSS nch l=0.04u w=0.4u
m9566 4974 4712 72205 VSS nch l=0.19u w=2.6u
m9567 4984 4977 VSS VSS nch l=0.04u w=0.8u
m9568 4993 4997 4990 VSS nch l=0.04u w=0.4u
m9569 4987 FOUT1PH270 VSS VSS nch l=0.04u w=0.4u
m9570 VSS 4977 4984 VSS nch l=0.04u w=0.8u
m9571 4995 4985 VSS VSS nch l=0.04u w=0.4u
m9572 72212 4712 4974 VSS nch l=0.19u w=2.6u
m9573 VSS FOUT1PH270 4987 VSS nch l=0.04u w=0.4u
m9574 4984 4977 VSS VSS nch l=0.04u w=0.8u
m9575 4997 5143 VSS VSS nch l=0.04u w=0.4u
m9576 VSS 4977 4984 VSS nch l=0.04u w=0.8u
m9577 VSS 4712 72212 VSS nch l=0.19u w=2.6u
m9578 4998 4995 4972 VSS nch l=0.04u w=0.4u
m9579 4999 4953 VSS VSS nch l=0.04u w=0.4u
m9580 4984 4977 VSS VSS nch l=0.04u w=0.8u
m9581 72218 4985 4998 VSS nch l=0.04u w=0.12u
m9582 72219 4712 VSS VSS nch l=0.19u w=2.6u
m9583 4989 4708 4984 VSS nch l=0.04u w=0.8u
m9584 VSS 5018 4993 VSS nch l=0.04u w=0.4u
m9585 VSS 5019 72218 VSS nch l=0.04u w=0.12u
m9586 4984 4708 4989 VSS nch l=0.04u w=0.8u
m9587 5019 4998 VSS VSS nch l=0.04u w=0.4u
m9588 4974 4712 72219 VSS nch l=0.19u w=2.6u
m9589 4989 4708 4984 VSS nch l=0.04u w=0.8u
m9590 VSS 5021 5017 VSS nch l=0.04u w=0.4u
m9591 72222 5023 5018 VSS nch l=0.04u w=0.8u
m9592 72227 4712 4974 VSS nch l=0.19u w=2.6u
m9593 VSS 4959 72222 VSS nch l=0.04u w=0.8u
m9594 5022 4985 5019 VSS nch l=0.04u w=0.4u
m9595 72228 5039 5021 VSS nch l=0.04u w=0.8u
m9596 VSS 5037 5016 VSS nch l=0.04u w=0.4u
m9597 5024 4989 VSS VSS nch l=0.04u w=0.4u
m9598 72229 4995 5022 VSS nch l=0.04u w=0.12u
m9599 VSS 4712 72227 VSS nch l=0.19u w=2.6u
m9600 VSS 4999 72228 VSS nch l=0.04u w=0.8u
m9601 VSS 5045 5023 VSS nch l=0.04u w=0.4u
m9602 VSS 5042 72229 VSS nch l=0.04u w=0.12u
m9603 72234 4712 VSS VSS nch l=0.19u w=2.6u
m9604 72235 4993 VSS VSS nch l=0.04u w=0.12u
m9605 VSS 2426 5037 VSS nch l=0.04u w=0.4u
m9606 5042 5022 VSS VSS nch l=0.04u w=0.4u
m9607 5041 5024 5038 VSS nch l=0.04u w=0.4u
m9608 5045 5088 72235 VSS nch l=0.04u w=0.12u
m9609 VSS 5049 5039 VSS nch l=0.04u w=0.4u
m9610 5044 5037 VSS VSS nch l=0.04u w=0.4u
m9611 72236 4989 5041 VSS nch l=0.04u w=0.12u
m9612 4974 4712 72234 VSS nch l=0.19u w=2.6u
m9613 5046 5143 5045 VSS nch l=0.04u w=0.4u
m9614 72237 5017 VSS VSS nch l=0.04u w=0.12u
m9615 VSS 5051 72236 VSS nch l=0.04u w=0.12u
m9616 5047 4863 VSS VSS nch l=0.04u w=0.4u
m9617 72238 4712 4974 VSS nch l=0.19u w=2.6u
m9618 5049 5094 72237 VSS nch l=0.04u w=0.12u
m9619 5050 5044 VSS VSS nch l=0.04u w=0.4u
m9620 5051 5041 VSS VSS nch l=0.04u w=0.4u
m9621 5064 5248 5049 VSS nch l=0.04u w=0.4u
m9622 72242 5069 5046 VSS nch l=0.04u w=0.8u
m9623 VSS 4712 72238 VSS nch l=0.19u w=2.6u
m9624 72243 4863 VSS VSS nch l=0.04u w=0.8u
m9625 VSS 4959 72242 VSS nch l=0.04u w=0.8u
m9626 5066 4989 5051 VSS nch l=0.04u w=0.4u
m9627 5065 5042 72243 VSS nch l=0.04u w=0.8u
m9628 VSS VSS VSS VSS nch l=0.19u w=2.6u
m9629 72247 5046 VSS VSS nch l=0.04u w=0.24u
m9630 72248 5085 5064 VSS nch l=0.04u w=0.8u
m9631 72249 5024 5066 VSS nch l=0.04u w=0.12u
m9632 5069 5143 72247 VSS nch l=0.04u w=0.24u
m9633 VSS 4999 72248 VSS nch l=0.04u w=0.8u
m9634 VSS 5071 72249 VSS nch l=0.04u w=0.12u
m9635 72250 5047 VSS VSS nch l=0.04u w=0.8u
m9636 4959 5088 5069 VSS nch l=0.04u w=0.4u
m9637 72251 5064 VSS VSS nch l=0.04u w=0.24u
m9638 5071 5066 VSS VSS nch l=0.04u w=0.4u
m9639 5070 4935 72250 VSS nch l=0.04u w=0.8u
m9640 5085 5248 72251 VSS nch l=0.04u w=0.24u
m9641 5087 5094 5085 VSS nch l=0.04u w=0.4u
m9642 5088 5143 VSS VSS nch l=0.04u w=0.4u
m9643 5089 4989 VSS VSS nch l=0.04u w=0.4u
m9644 72259 5070 VSS VSS nch l=0.04u w=0.8u
m9645 5090 5065 72259 VSS nch l=0.04u w=0.8u
m9646 5094 5248 VSS VSS nch l=0.04u w=0.4u
m9647 FOUT2 5132 VSS VSS nch l=0.04u w=0.4u
m9648 5096 5089 5071 VSS nch l=0.04u w=0.4u
m9649 72265 5065 5090 VSS nch l=0.04u w=0.8u
m9650 VSS 5132 FOUT2 VSS nch l=0.04u w=0.4u
m9651 72271 4989 5096 VSS nch l=0.04u w=0.12u
m9652 VSS 5070 72265 VSS nch l=0.04u w=0.8u
m9653 FOUT2 5132 VSS VSS nch l=0.04u w=0.4u
m9654 VSS 5111 72271 VSS nch l=0.04u w=0.12u
m9655 VSS 5112 5087 VSS nch l=0.04u w=0.4u
m9656 VSS 5132 FOUT2 VSS nch l=0.04u w=0.4u
m9657 5111 5096 VSS VSS nch l=0.04u w=0.4u
m9658 VSS 4858 5110 VSS nch l=0.04u w=0.8u
m9659 FOUT2 5132 VSS VSS nch l=0.04u w=0.4u
m9660 72273 5117 5112 VSS nch l=0.04u w=0.8u
m9661 5110 4858 VSS VSS nch l=0.04u w=0.8u
m9662 VSS 5132 FOUT2 VSS nch l=0.04u w=0.4u
m9663 5115 4989 5111 VSS nch l=0.04u w=0.4u
m9664 VSS 4999 72273 VSS nch l=0.04u w=0.8u
m9665 5113 5527 5110 VSS nch l=0.04u w=0.8u
m9666 FOUT2 5132 VSS VSS nch l=0.04u w=0.4u
m9667 72278 5089 5115 VSS nch l=0.04u w=0.12u
m9668 VSS 5132 FOUT2 VSS nch l=0.04u w=0.4u
m9669 VSS 5133 72278 VSS nch l=0.04u w=0.12u
m9670 VSS 5135 5117 VSS nch l=0.04u w=0.4u
m9671 5130 5113 VSS VSS nch l=0.04u w=0.4u
m9672 5133 5115 VSS VSS nch l=0.04u w=0.4u
m9673 72282 5087 VSS VSS nch l=0.04u w=0.12u
m9674 VSS 5137 5116 VSS nch l=0.04u w=0.4u
m9675 5134 5162 5132 VSS nch l=0.04u w=0.8u
m9676 5135 5182 72282 VSS nch l=0.04u w=0.12u
m9677 5136 5130 5090 VSS nch l=0.04u w=0.4u
m9678 VSS 4962 5134 VSS nch l=0.04u w=0.8u
m9679 5138 5248 5135 VSS nch l=0.04u w=0.4u
m9680 72287 5113 5136 VSS nch l=0.04u w=0.12u
m9681 VSS 2427 5137 VSS nch l=0.04u w=0.4u
m9682 5134 4962 VSS VSS nch l=0.04u w=0.8u
m9683 5140 4989 VSS VSS nch l=0.04u w=0.4u
m9684 VSS 5156 72287 VSS nch l=0.04u w=0.12u
m9685 5142 5137 VSS VSS nch l=0.04u w=0.4u
m9686 72289 5163 5138 VSS nch l=0.04u w=0.8u
m9687 5156 5136 VSS VSS nch l=0.04u w=0.4u
m9688 VSS 5160 5143 VSS nch l=0.04u w=0.4u
m9689 5157 5140 5133 VSS nch l=0.04u w=0.4u
m9690 VSS 4999 72289 VSS nch l=0.04u w=0.8u
m9691 5159 5142 VSS VSS nch l=0.04u w=0.4u
m9692 5160 5162 VSS VSS nch l=0.04u w=0.4u
m9693 72290 4989 5157 VSS nch l=0.04u w=0.12u
m9694 72291 5138 VSS VSS nch l=0.04u w=0.24u
m9695 5161 5113 5156 VSS nch l=0.04u w=0.4u
m9696 VSS 5164 72290 VSS nch l=0.04u w=0.12u
m9697 5163 5248 72291 VSS nch l=0.04u w=0.24u
m9698 72296 5130 5161 VSS nch l=0.04u w=0.12u
m9699 72297 5204 5162 VSS nch l=0.04u w=0.8u
m9700 5164 5157 VSS VSS nch l=0.04u w=0.4u
m9701 4999 5182 5163 VSS nch l=0.04u w=0.4u
m9702 VSS 5177 72296 VSS nch l=0.04u w=0.12u
m9703 VSS 5180 72297 VSS nch l=0.04u w=0.8u
m9704 5177 5161 VSS VSS nch l=0.04u w=0.4u
m9705 5181 4989 5164 VSS nch l=0.04u w=0.4u
m9706 5182 5248 VSS VSS nch l=0.04u w=0.4u
m9707 VSS 5179 5179 VSS nch l=0.04u w=0.8u
m9708 72304 5140 5181 VSS nch l=0.04u w=0.12u
m9709 VSS 5189 72304 VSS nch l=0.04u w=0.12u
m9710 5185 5186 VSS VSS nch l=0.04u w=0.8u
m9711 FOUT1PH180 5226 VSS VSS nch l=0.04u w=0.4u
m9712 5188 5177 VSS VSS nch l=0.04u w=0.4u
m9713 VSS 5204 5184 VSS nch l=0.04u w=0.4u
m9714 5189 5181 VSS VSS nch l=0.04u w=0.4u
m9715 VSS 5226 FOUT1PH180 VSS nch l=0.04u w=0.4u
m9716 FOUT1PH180 5226 VSS VSS nch l=0.04u w=0.4u
m9717 72315 4876 VSS VSS nch l=0.04u w=0.8u
m9718 VSS 5226 FOUT1PH180 VSS nch l=0.04u w=0.4u
m9719 72320 5188 72315 VSS nch l=0.04u w=0.8u
m9720 VSS 5210 5204 VSS nch l=0.04u w=0.4u
m9721 FOUT1PH180 5226 VSS VSS nch l=0.04u w=0.4u
m9722 5203 5042 72320 VSS nch l=0.04u w=0.8u
m9723 5207 4989 VSS VSS nch l=0.04u w=0.4u
m9724 72323 5204 VSS VSS nch l=0.04u w=0.12u
m9725 VSS 5226 FOUT1PH180 VSS nch l=0.04u w=0.4u
m9726 5210 5257 72323 VSS nch l=0.04u w=0.12u
m9727 FOUT1PH180 5226 VSS VSS nch l=0.04u w=0.4u
m9728 VSS 5206 5208 VSS nch l=0.04u w=0.4u
m9729 VSS POSTDIV2[0] 5209 VSS nch l=0.04u w=0.8u
m9730 5211 5207 5189 VSS nch l=0.04u w=0.4u
m9731 5213 5277 5210 VSS nch l=0.04u w=0.4u
m9732 VSS 5226 FOUT1PH180 VSS nch l=0.04u w=0.4u
m9733 5209 POSTDIV2[0] VSS VSS nch l=0.04u w=0.8u
m9734 72332 4989 5211 VSS nch l=0.04u w=0.12u
m9735 5212 5188 5209 VSS nch l=0.04u w=0.62u
m9736 5227 5230 VSS VSS nch l=0.04u w=0.4u
m9737 VSS 5229 72332 VSS nch l=0.04u w=0.12u
m9738 VSS 5233 5213 VSS nch l=0.04u w=0.4u
m9739 5228 5343 5226 VSS nch l=0.04u w=0.8u
m9740 5229 5211 VSS VSS nch l=0.04u w=0.4u
m9741 72336 5213 VSS VSS nch l=0.04u w=0.12u
m9742 VSS 5017 5228 VSS nch l=0.04u w=0.8u
m9743 72337 5203 VSS VSS nch l=0.04u w=0.8u
m9744 5233 5277 72336 VSS nch l=0.04u w=0.12u
m9745 5228 5017 VSS VSS nch l=0.04u w=0.8u
m9746 5235 4989 5229 VSS nch l=0.04u w=0.4u
m9747 72346 5212 72337 VSS nch l=0.04u w=0.8u
m9748 72349 5208 5232 VSS nch l=0.04u w=0.8u
m9749 5184 5257 5233 VSS nch l=0.04u w=0.4u
m9750 72350 5207 5235 VSS nch l=0.04u w=0.12u
m9751 4935 5439 72346 VSS nch l=0.04u w=0.8u
m9752 VSS 5271 72349 VSS nch l=0.04u w=0.8u
m9753 VSS 5253 5248 VSS nch l=0.04u w=0.4u
m9754 VSS 5254 72350 VSS nch l=0.04u w=0.12u
m9755 5253 5343 VSS VSS nch l=0.04u w=0.4u
m9756 5254 5235 VSS VSS nch l=0.04u w=0.4u
m9757 72354 5203 VSS VSS nch l=0.04u w=0.8u
m9758 5255 5257 5252 VSS nch l=0.04u w=0.4u
m9759 72359 5212 72354 VSS nch l=0.04u w=0.8u
m9760 72360 5277 5255 VSS nch l=0.04u w=0.12u
m9761 VSS 5251 5256 VSS nch l=0.04u w=0.4u
m9762 5257 5277 VSS VSS nch l=0.04u w=0.4u
m9763 72361 5189 VSS VSS nch l=0.04u w=0.8u
m9764 4935 5439 72359 VSS nch l=0.04u w=0.8u
m9765 VSS 5270 72360 VSS nch l=0.04u w=0.12u
m9766 VSS 5277 5257 VSS nch l=0.04u w=0.4u
m9767 5038 5254 72361 VSS nch l=0.04u w=0.8u
m9768 5270 5255 VSS VSS nch l=0.04u w=0.4u
m9769 5271 5274 VSS VSS nch l=0.04u w=0.4u
m9770 5257 5277 VSS VSS nch l=0.04u w=0.4u
m9771 72366 5254 5038 VSS nch l=0.04u w=0.8u
m9772 5272 4858 VSS VSS nch l=0.04u w=0.4u
m9773 VSS 5277 5257 VSS nch l=0.04u w=0.4u
m9774 VSS 5189 72366 VSS nch l=0.04u w=0.8u
m9775 5275 5277 5270 VSS nch l=0.04u w=0.4u
m9776 72375 5257 5275 VSS nch l=0.04u w=0.12u
m9777 72376 4858 VSS VSS nch l=0.04u w=0.8u
m9778 5277 FOUT1PH180 VSS VSS nch l=0.04u w=0.4u
m9779 5278 5229 VSS VSS nch l=0.04u w=0.4u
m9780 VSS 5291 72375 VSS nch l=0.04u w=0.12u
m9781 5276 5177 72376 VSS nch l=0.04u w=0.8u
m9782 VSS FOUT1PH180 5277 VSS nch l=0.04u w=0.4u
m9783 5291 5275 VSS VSS nch l=0.04u w=0.4u
m9784 5277 FOUT1PH180 VSS VSS nch l=0.04u w=0.4u
m9785 72391 4977 VSS VSS nch l=0.04u w=0.8u
m9786 72392 5272 VSS VSS nch l=0.04u w=0.8u
m9787 VSS FOUT1PH180 5277 VSS nch l=0.04u w=0.4u
m9788 72395 5278 72391 VSS nch l=0.04u w=0.8u
m9789 5294 5291 VSS VSS nch l=0.04u w=0.4u
m9790 5293 4935 72392 VSS nch l=0.04u w=0.8u
m9791 5292 5254 72395 VSS nch l=0.04u w=0.8u
m9792 5252 5204 5294 VSS nch l=0.04u w=0.4u
m9793 5295 FOUTPOSTDIV VSS VSS nch l=0.04u w=0.4u
m9794 5204 5294 5252 VSS nch l=0.04u w=0.4u
m9795 72402 5293 VSS VSS nch l=0.04u w=0.8u
m9796 VSS 4956 5296 VSS nch l=0.04u w=0.8u
m9797 5297 5276 72402 VSS nch l=0.04u w=0.8u
m9798 5311 5295 VSS VSS nch l=0.04u w=0.4u
m9799 5296 4956 VSS VSS nch l=0.04u w=0.8u
m9800 72408 5276 5297 VSS nch l=0.04u w=0.8u
m9801 VSS 5295 5311 VSS nch l=0.04u w=0.4u
m9802 5310 4708 5296 VSS nch l=0.04u w=0.8u
m9803 VSS 5293 72408 VSS nch l=0.04u w=0.8u
m9804 5317 5317 VSS VSS nch l=0.04u w=0.8u
m9805 5320 5311 5319 VSS nch l=0.04u w=0.4u
m9806 5321 5310 VSS VSS nch l=0.04u w=0.4u
m9807 5323 5323 VSS VSS nch l=0.04u w=0.8u
m9808 72409 5318 VSS VSS nch l=0.04u w=0.8u
m9809 72414 5295 5320 VSS nch l=0.04u w=0.12u
m9810 5324 5291 72409 VSS nch l=0.04u w=0.8u
m9811 VSS 5343 72414 VSS nch l=0.04u w=0.12u
m9812 5340 5321 5337 VSS nch l=0.04u w=0.4u
m9813 VSS 5322 5338 VSS nch l=0.04u w=0.8u
m9814 5343 5320 VSS VSS nch l=0.04u w=0.4u
m9815 72415 5310 5340 VSS nch l=0.04u w=0.12u
m9816 5338 5322 VSS VSS nch l=0.04u w=0.8u
m9817 VSS 5324 5342 VSS nch l=0.04u w=0.4u
m9818 VSS 5362 72415 VSS nch l=0.04u w=0.12u
m9819 5341 5527 5338 VSS nch l=0.04u w=0.8u
m9820 5361 5342 VSS VSS nch l=0.04u w=0.4u
m9821 5362 5340 VSS VSS nch l=0.04u w=0.4u
m9822 5363 5343 VSS VSS nch l=0.04u w=0.4u
m9823 VSS 5343 5363 VSS nch l=0.04u w=0.4u
m9824 5377 5341 VSS VSS nch l=0.04u w=0.4u
m9825 VSS 5676 5364 VSS nch l=0.04u w=0.8u
m9826 5379 5310 5362 VSS nch l=0.04u w=0.4u
m9827 5364 5676 VSS VSS nch l=0.04u w=0.8u
m9828 72422 5321 5379 VSS nch l=0.04u w=0.12u
m9829 5392 5343 VSS VSS nch l=0.04u w=0.4u
m9830 5378 5324 5364 VSS nch l=0.04u w=0.8u
m9831 5393 5377 5297 VSS nch l=0.04u w=0.4u
m9832 VSS 5394 72422 VSS nch l=0.04u w=0.12u
m9833 72431 5341 5393 VSS nch l=0.04u w=0.12u
m9834 5394 5379 VSS VSS nch l=0.04u w=0.4u
m9835 VSS 5409 72431 VSS nch l=0.04u w=0.12u
m9836 FOUT4 5378 VSS VSS nch l=0.04u w=0.4u
m9837 5396 5295 5392 VSS nch l=0.04u w=0.4u
m9838 5409 5393 VSS VSS nch l=0.04u w=0.4u
m9839 VSS 5378 FOUT4 VSS nch l=0.04u w=0.4u
m9840 72446 5311 5396 VSS nch l=0.04u w=0.12u
m9841 FOUT4 5378 VSS VSS nch l=0.04u w=0.4u
m9842 VSS 5424 72446 VSS nch l=0.04u w=0.12u
m9843 5410 5310 VSS VSS nch l=0.04u w=0.4u
m9844 VSS 5378 FOUT4 VSS nch l=0.04u w=0.4u
m9845 5423 5341 5409 VSS nch l=0.04u w=0.4u
m9846 5424 5396 VSS VSS nch l=0.04u w=0.4u
m9847 FOUT4 5378 VSS VSS nch l=0.04u w=0.4u
m9848 72451 5377 5423 VSS nch l=0.04u w=0.12u
m9849 5425 5410 5394 VSS nch l=0.04u w=0.4u
m9850 VSS 5378 FOUT4 VSS nch l=0.04u w=0.4u
m9851 VSS 5439 72451 VSS nch l=0.04u w=0.12u
m9852 5426 5424 VSS VSS nch l=0.04u w=0.4u
m9853 72478 5310 5425 VSS nch l=0.04u w=0.12u
m9854 FOUT4 5378 VSS VSS nch l=0.04u w=0.4u
m9855 5439 5423 VSS VSS nch l=0.04u w=0.4u
m9856 VSS 5424 5426 VSS nch l=0.04u w=0.4u
m9857 VSS 5440 72478 VSS nch l=0.04u w=0.12u
m9858 VSS 5378 FOUT4 VSS nch l=0.04u w=0.4u
m9859 5440 5425 VSS VSS nch l=0.04u w=0.4u
m9860 5455 5424 VSS VSS nch l=0.04u w=0.4u
m9861 VSS POSTDIV2[0] 5441 VSS nch l=0.04u w=0.8u
m9862 VSS 5361 5454 VSS nch l=0.04u w=0.4u
m9863 5441 POSTDIV2[0] VSS VSS nch l=0.04u w=0.8u
m9864 5457 5310 5440 VSS nch l=0.04u w=0.4u
m9865 5319 5455 VSS VSS nch l=0.04u w=0.4u
m9866 5456 5409 5441 VSS nch l=0.04u w=0.62u
m9867 72512 5410 5457 VSS nch l=0.04u w=0.12u
m9868 5471 5454 5458 VSS nch l=0.04u w=0.4u
m9869 VSS 5473 72512 VSS nch l=0.04u w=0.12u
m9870 72514 5361 5471 VSS nch l=0.04u w=0.24u
m9871 5472 FOUT1PH90 VSS VSS nch l=0.04u w=0.4u
m9872 5473 5457 VSS VSS nch l=0.04u w=0.4u
m9873 VSS 5487 72514 VSS nch l=0.04u w=0.24u
m9874 72527 5456 VSS VSS nch l=0.04u w=0.8u
m9875 VSS FOUT1PH90 5472 VSS nch l=0.04u w=0.4u
m9876 72539 5458 VSS VSS nch l=0.04u w=0.8u
m9877 5486 5439 72527 VSS nch l=0.04u w=0.8u
m9878 5472 FOUT1PH90 VSS VSS nch l=0.04u w=0.4u
m9879 5487 5471 72539 VSS nch l=0.04u w=0.8u
m9880 VSS FOUT1PH90 5472 VSS nch l=0.04u w=0.4u
m9881 5503 5310 VSS VSS nch l=0.04u w=0.4u
m9882 5339 5814 5488 VSS nch l=0.25u w=0.65u
m9883 5339 5814 5488 VSS nch l=0.25u w=0.65u
m9884 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9885 5504 5486 VSS VSS nch l=0.04u w=0.4u
m9886 72551 5784 VSS VSS nch l=0.25u w=0.5u
m9887 72552 5732 VSS VSS nch l=0.25u w=0.5u
m9888 5508 5361 5487 VSS nch l=0.04u w=0.4u
m9889 VSS 5486 5504 VSS nch l=0.04u w=0.4u
m9890 VSS 5426 5505 VSS nch l=0.04u w=0.4u
m9891 5488 5814 5339 VSS nch l=0.25u w=0.65u
m9892 5488 5814 5339 VSS nch l=0.25u w=0.65u
m9893 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9894 5511 5510 5507 VSS nch l=0.13u w=1.3u
m9895 72557 5454 5508 VSS nch l=0.04u w=0.12u
m9896 5512 5503 5473 VSS nch l=0.04u w=0.4u
m9897 72558 5784 72551 VSS nch l=0.25u w=0.5u
m9898 72559 5732 72552 VSS nch l=0.25u w=0.5u
m9899 5525 5505 VSS VSS nch l=0.04u w=0.4u
m9900 VSS 5564 72557 VSS nch l=0.04u w=0.12u
m9901 72565 5310 5512 VSS nch l=0.04u w=0.12u
m9902 5527 5549 VSS VSS nch l=0.04u w=0.4u
m9903 5507 5510 5511 VSS nch l=0.13u w=1.3u
m9904 5528 5814 5509 VSS nch l=0.25u w=0.65u
m9905 5339 5814 5488 VSS nch l=0.25u w=0.65u
m9906 5339 5814 5488 VSS nch l=0.25u w=0.65u
m9907 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9908 5531 5508 VSS VSS nch l=0.04u w=0.4u
m9909 72567 5784 72558 VSS nch l=0.25u w=0.5u
m9910 72568 5732 72559 VSS nch l=0.25u w=0.5u
m9911 VSS 5534 72565 VSS nch l=0.04u w=0.12u
m9912 VSS 5549 5527 VSS nch l=0.04u w=0.4u
m9913 5526 5532 5507 VSS nch l=0.13u w=1.3u
m9914 VSS 5794 5530 VSS nch l=0.04u w=0.8u
m9915 5509 5814 5528 VSS nch l=0.25u w=0.65u
m9916 5534 5512 VSS VSS nch l=0.04u w=0.4u
m9917 5488 5814 5339 VSS nch l=0.25u w=0.65u
m9918 5488 5814 5339 VSS nch l=0.25u w=0.65u
m9919 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9920 5530 5794 VSS VSS nch l=0.04u w=0.8u
m9921 5507 5532 5526 VSS nch l=0.13u w=1.3u
m9922 5547 5784 72567 VSS nch l=0.25u w=0.5u
m9923 5509 5732 72568 VSS nch l=0.25u w=0.5u
m9924 72574 5458 VSS VSS nch l=0.04u w=0.8u
m9925 72580 4710 VSS VSS nch l=0.04u w=0.8u
m9926 5533 5426 5530 VSS nch l=0.04u w=0.8u
m9927 5511 5510 5507 VSS nch l=0.13u w=1.3u
m9928 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9929 5548 5531 72574 VSS nch l=0.04u w=0.8u
m9930 5550 5310 5534 VSS nch l=0.04u w=0.4u
m9931 72582 5767 72580 VSS nch l=0.04u w=0.8u
m9932 72584 5784 5547 VSS nch l=0.25u w=0.5u
m9933 72585 5732 5509 VSS nch l=0.25u w=0.5u
m9934 72586 5503 5550 VSS nch l=0.04u w=0.12u
m9935 5507 5510 5511 VSS nch l=0.13u w=1.3u
m9936 5549 5580 72582 VSS nch l=0.04u w=0.8u
m9937 5532 5814 5547 VSS nch l=0.25u w=0.65u
m9938 72587 5784 VSS VSS nch l=0.25u w=0.5u
m9939 72588 5784 VSS VSS nch l=0.25u w=0.5u
m9940 FOUT1PH90 5533 VSS VSS nch l=0.04u w=0.4u
m9941 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9942 VSS 5566 72586 VSS nch l=0.04u w=0.12u
m9943 5564 5548 VSS VSS nch l=0.04u w=0.4u
m9944 5526 5532 5507 VSS nch l=0.13u w=1.3u
m9945 72594 5784 72584 VSS nch l=0.25u w=0.5u
m9946 72595 5732 72585 VSS nch l=0.25u w=0.5u
m9947 VSS 5533 FOUT1PH90 VSS nch l=0.04u w=0.4u
m9948 5566 5550 VSS VSS nch l=0.04u w=0.4u
m9949 5547 5814 5532 VSS nch l=0.25u w=0.65u
m9950 72601 5784 72587 VSS nch l=0.25u w=0.5u
m9951 72602 5784 72588 VSS nch l=0.25u w=0.5u
m9952 VSS 4715 5565 VSS nch l=0.04u w=0.8u
m9953 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9954 FOUT1PH90 5533 VSS VSS nch l=0.04u w=0.4u
m9955 5507 5532 5526 VSS nch l=0.13u w=1.3u
m9956 72606 5784 72594 VSS nch l=0.25u w=0.5u
m9957 72607 5732 72595 VSS nch l=0.25u w=0.5u
m9958 5565 4715 VSS VSS nch l=0.04u w=0.8u
m9959 VSS 5361 5579 VSS nch l=0.04u w=0.4u
m9960 VSS 5533 FOUT1PH90 VSS nch l=0.04u w=0.4u
m9961 5511 5510 5507 VSS nch l=0.13u w=1.3u
m9962 72612 5784 72601 VSS nch l=0.25u w=0.5u
m9963 72613 5784 72602 VSS nch l=0.25u w=0.5u
m9964 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9965 VSS POSTDIV1[0] 5581 VSS nch l=0.04u w=0.8u
m9966 5580 4708 5565 VSS nch l=0.04u w=0.62u
m9967 FOUT1PH90 5533 VSS VSS nch l=0.04u w=0.4u
m9968 5507 5510 5511 VSS nch l=0.13u w=1.3u
m9969 VSS 5784 72606 VSS nch l=0.25u w=0.5u
m9970 VSS 5732 72607 VSS nch l=0.25u w=0.5u
m9971 5581 POSTDIV1[0] VSS VSS nch l=0.04u w=0.8u
m9972 5596 5579 5564 VSS nch l=0.04u w=0.4u
m9973 VSS 5533 FOUT1PH90 VSS nch l=0.04u w=0.4u
m9974 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9975 5488 5784 72612 VSS nch l=0.25u w=0.5u
m9976 5488 5784 72613 VSS nch l=0.25u w=0.5u
m9977 5594 5534 5581 VSS nch l=0.04u w=0.62u
m9978 5526 5532 5507 VSS nch l=0.13u w=1.3u
m9979 72616 5361 5596 VSS nch l=0.04u w=0.24u
m9980 FOUT1PH90 5533 VSS VSS nch l=0.04u w=0.4u
m9981 5597 4860 VSS VSS nch l=0.04u w=0.4u
m9982 72619 5784 VSS VSS nch l=0.25u w=0.5u
m9983 72620 5784 VSS VSS nch l=0.25u w=0.5u
m9984 5532 4 VDDREF VSS nch l=0.1u w=1.3u
m9985 VSS 5612 72616 VSS nch l=0.04u w=0.24u
m9986 VSS 5533 FOUT1PH90 VSS nch l=0.04u w=0.4u
m9987 5507 5532 5526 VSS nch l=0.13u w=1.3u
m9988 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m9989 72623 5784 5488 VSS nch l=0.25u w=0.5u
m9990 72624 5784 5488 VSS nch l=0.25u w=0.5u
m9991 VDDREF 4 5532 VSS nch l=0.1u w=1.3u
m9992 72627 4956 VSS VSS nch l=0.04u w=0.8u
m9993 72628 5458 VSS VSS nch l=0.04u w=0.8u
m9994 72630 4860 VSS VSS nch l=0.04u w=0.8u
m9995 5511 5510 5507 VSS nch l=0.13u w=1.3u
m9996 72631 5784 72619 VSS nch l=0.25u w=0.5u
m9997 72632 5784 72620 VSS nch l=0.25u w=0.5u
m9998 5532 4 VDDREF VSS nch l=0.1u w=1.3u
m9999 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10000 72637 5594 72627 VSS nch l=0.04u w=0.8u
m10001 5612 5596 72628 VSS nch l=0.04u w=0.8u
m10002 VSS 5525 5613 VSS nch l=0.04u w=0.4u
m10003 72639 5784 72623 VSS nch l=0.25u w=0.5u
m10004 72640 5784 72624 VSS nch l=0.25u w=0.5u
m10005 5614 4707 72630 VSS nch l=0.04u w=0.8u
m10006 5507 5510 5511 VSS nch l=0.13u w=1.3u
m10007 VDDREF 4 5532 VSS nch l=0.1u w=1.3u
m10008 5611 5566 72637 VSS nch l=0.04u w=0.8u
m10009 72644 5784 72631 VSS nch l=0.25u w=0.5u
m10010 72645 5784 72632 VSS nch l=0.25u w=0.5u
m10011 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10012 5526 5532 5507 VSS nch l=0.13u w=1.3u
m10013 5532 4 VDDREF VSS nch l=0.1u w=1.3u
m10014 5628 5361 5612 VSS nch l=0.04u w=0.4u
m10015 72646 5784 72639 VSS nch l=0.25u w=0.5u
m10016 72647 5784 72640 VSS nch l=0.25u w=0.5u
m10017 5629 5613 5627 VSS nch l=0.04u w=0.4u
m10018 72655 5597 VSS VSS nch l=0.04u w=0.8u
m10019 72656 5566 5337 VSS nch l=0.04u w=0.8u
m10020 72657 5579 5628 VSS nch l=0.04u w=0.12u
m10021 5507 5532 5526 VSS nch l=0.13u w=1.3u
m10022 5507 5784 72644 VSS nch l=0.25u w=0.5u
m10023 5507 5784 72645 VSS nch l=0.25u w=0.5u
m10024 VDDREF 4 5532 VSS nch l=0.1u w=1.3u
m10025 72658 5525 5629 VSS nch l=0.04u w=0.24u
m10026 5630 5504 72655 VSS nch l=0.04u w=0.8u
m10027 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10028 VSS 5784 72646 VSS nch l=0.25u w=0.5u
m10029 VSS 5784 72647 VSS nch l=0.25u w=0.5u
m10030 72661 5660 72656 VSS nch l=0.04u w=0.8u
m10031 VSS 5676 72657 VSS nch l=0.04u w=0.12u
m10032 VSS 5657 72658 VSS nch l=0.04u w=0.24u
m10033 5510 5015 VDDREF VSS nch l=0.1u w=1.3u
m10034 5526 5532 5507 VSS nch l=0.13u w=1.3u
m10035 72669 5784 5507 VSS nch l=0.25u w=0.5u
m10036 72670 5784 5507 VSS nch l=0.25u w=0.5u
m10037 VSS 5693 72661 VSS nch l=0.04u w=0.8u
m10038 5644 5628 VSS VSS nch l=0.04u w=0.4u
m10039 72671 5627 VSS VSS nch l=0.04u w=0.8u
m10040 VDDREF 5015 5510 VSS nch l=0.1u w=1.3u
m10041 72672 5630 VSS VSS nch l=0.04u w=0.8u
m10042 5507 5532 5526 VSS nch l=0.13u w=1.3u
m10043 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10044 72673 5784 VSS VSS nch l=0.25u w=0.5u
m10045 72674 5784 VSS VSS nch l=0.25u w=0.5u
m10046 5657 5629 72671 VSS nch l=0.04u w=0.8u
m10047 5510 5015 VDDREF VSS nch l=0.1u w=1.3u
m10048 5658 5614 72672 VSS nch l=0.04u w=0.8u
m10049 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10050 72682 5784 72669 VSS nch l=0.25u w=0.5u
m10051 72683 5784 72670 VSS nch l=0.25u w=0.5u
m10052 5511 5510 5507 VSS nch l=0.13u w=1.3u
m10053 72684 5458 VSS VSS nch l=0.04u w=0.8u
m10054 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10055 5662 5690 5660 VSS nch l=0.04u w=0.62u
m10056 72688 5614 5658 VSS nch l=0.04u w=0.8u
m10057 VDDREF 5015 5510 VSS nch l=0.1u w=1.3u
m10058 72689 5784 72673 VSS nch l=0.25u w=0.5u
m10059 72690 5784 72674 VSS nch l=0.25u w=0.5u
m10060 5507 5510 5511 VSS nch l=0.13u w=1.3u
m10061 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10062 5661 5644 72684 VSS nch l=0.04u w=0.8u
m10063 5675 5525 5657 VSS nch l=0.04u w=0.4u
m10064 VSS POSTDIV1[0] 5662 VSS nch l=0.04u w=0.8u
m10065 VSS 5630 72688 VSS nch l=0.04u w=0.8u
m10066 5510 5015 VDDREF VSS nch l=0.1u w=1.3u
m10067 72697 5784 72682 VSS nch l=0.25u w=0.5u
m10068 72698 5784 72683 VSS nch l=0.25u w=0.5u
m10069 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10070 72699 5613 5675 VSS nch l=0.04u w=0.12u
m10071 5662 POSTDIV1[0] VSS VSS nch l=0.04u w=0.8u
m10072 5526 5532 5507 VSS nch l=0.13u w=1.3u
m10073 72704 5784 72689 VSS nch l=0.25u w=0.5u
m10074 72705 5784 72690 VSS nch l=0.25u w=0.5u
m10075 VDDREF 5015 5510 VSS nch l=0.1u w=1.3u
m10076 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10077 5676 5661 VSS VSS nch l=0.04u w=0.4u
m10078 VSS 5724 72699 VSS nch l=0.04u w=0.12u
m10079 5689 4711 VSS VSS nch l=0.04u w=0.4u
m10080 VSS 5784 72697 VSS nch l=0.25u w=0.5u
m10081 VSS 5784 72698 VSS nch l=0.25u w=0.5u
m10082 5507 5532 5526 VSS nch l=0.13u w=1.3u
m10083 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10084 5691 5675 VSS VSS nch l=0.04u w=0.4u
m10085 5488 5784 72704 VSS nch l=0.25u w=0.5u
m10086 5488 5784 72705 VSS nch l=0.25u w=0.5u
m10087 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10088 VSS 5473 5690 VSS nch l=0.04u w=0.4u
m10089 5511 5510 5507 VSS nch l=0.13u w=1.3u
m10090 72720 5784 VSS VSS nch l=0.25u w=0.5u
m10091 72721 5732 VSS VSS nch l=0.25u w=0.5u
m10092 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10093 72722 4711 VSS VSS nch l=0.04u w=0.8u
m10094 5507 5510 5511 VSS nch l=0.13u w=1.3u
m10095 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10096 72724 5784 5488 VSS nch l=0.25u w=0.5u
m10097 72725 5784 5488 VSS nch l=0.25u w=0.5u
m10098 72726 5627 VSS VSS nch l=0.04u w=0.8u
m10099 VSS 4953 5458 VSS nch l=0.04u w=0.4u
m10100 5692 5767 72722 VSS nch l=0.04u w=0.8u
m10101 72727 5394 5693 VSS nch l=0.04u w=0.8u
m10102 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10103 72729 5784 72720 VSS nch l=0.25u w=0.5u
m10104 72730 5732 72721 VSS nch l=0.25u w=0.5u
m10105 5706 5691 72726 VSS nch l=0.04u w=0.8u
m10106 5526 5532 5507 VSS nch l=0.13u w=1.3u
m10107 72731 5690 72727 VSS nch l=0.04u w=0.8u
m10108 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10109 72734 5784 72724 VSS nch l=0.25u w=0.5u
m10110 72735 5784 72725 VSS nch l=0.25u w=0.5u
m10111 5510 5814 5707 VSS nch l=0.25u w=0.65u
m10112 5507 5532 5526 VSS nch l=0.13u w=1.3u
m10113 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10114 VSS 4965 72731 VSS nch l=0.04u w=0.8u
m10115 72738 5689 VSS VSS nch l=0.04u w=0.8u
m10116 5722 5277 5708 VSS nch l=0.04u w=0.4u
m10117 72740 5784 72729 VSS nch l=0.25u w=0.5u
m10118 72741 5732 72730 VSS nch l=0.25u w=0.5u
m10119 5724 5706 VSS VSS nch l=0.04u w=0.4u
m10120 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10121 5721 5658 72738 VSS nch l=0.04u w=0.8u
m10122 72743 5257 5722 VSS nch l=0.04u w=0.12u
m10123 5511 5510 5507 VSS nch l=0.13u w=1.3u
m10124 72744 5784 72734 VSS nch l=0.25u w=0.5u
m10125 72745 5784 72735 VSS nch l=0.25u w=0.5u
m10126 5707 5814 5510 VSS nch l=0.25u w=0.65u
m10127 5015 5528 VSS VSS nch l=0.04u w=1.3u
m10128 72749 5292 VSS VSS nch l=0.04u w=0.8u
m10129 VSS 5731 72743 VSS nch l=0.04u w=0.12u
m10130 5707 5784 72740 VSS nch l=0.25u w=0.5u
m10131 5729 5732 72741 VSS nch l=0.25u w=0.5u
m10132 5507 5510 5511 VSS nch l=0.13u w=1.3u
m10133 VSS 5528 5015 VSS nch l=0.04u w=1.3u
m10134 72752 5611 72749 VSS nch l=0.04u w=0.8u
m10135 72753 5721 VSS VSS nch l=0.04u w=0.8u
m10136 5731 5722 VSS VSS nch l=0.04u w=0.4u
m10137 VSS 5525 5728 VSS nch l=0.04u w=0.4u
m10138 VSS 5784 72744 VSS nch l=0.25u w=0.5u
m10139 VSS 5784 72745 VSS nch l=0.25u w=0.5u
m10140 5526 5532 5507 VSS nch l=0.13u w=1.3u
m10141 72758 5784 5707 VSS nch l=0.25u w=0.5u
m10142 72759 5732 5729 VSS nch l=0.25u w=0.5u
m10143 5727 5798 72752 VSS nch l=0.04u w=0.8u
m10144 5730 5692 72753 VSS nch l=0.04u w=0.8u
m10145 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10146 5732 5814 5729 VSS nch l=0.25u w=0.65u
m10147 72761 5784 VSS VSS nch l=0.25u w=0.5u
m10148 72762 5784 VSS VSS nch l=0.25u w=0.5u
m10149 5507 5532 5526 VSS nch l=0.13u w=1.3u
m10150 72763 5692 5730 VSS nch l=0.04u w=0.8u
m10151 5746 5257 5731 VSS nch l=0.04u w=0.4u
m10152 5747 5728 5724 VSS nch l=0.04u w=0.4u
m10153 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10154 72765 5784 72758 VSS nch l=0.25u w=0.5u
m10155 72766 5732 72759 VSS nch l=0.25u w=0.5u
m10156 VSS 5721 72763 VSS nch l=0.04u w=0.8u
m10157 5748 5727 VSS VSS nch l=0.04u w=0.4u
m10158 72767 5277 5746 VSS nch l=0.04u w=0.12u
m10159 72768 5525 5747 VSS nch l=0.04u w=0.24u
m10160 5511 5510 5507 VSS nch l=0.13u w=1.3u
m10161 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10162 5729 5814 5732 VSS nch l=0.25u w=0.65u
m10163 72774 5784 72761 VSS nch l=0.25u w=0.5u
m10164 72775 5784 72762 VSS nch l=0.25u w=0.5u
m10165 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10166 VSS 5750 72767 VSS nch l=0.04u w=0.12u
m10167 VSS 5751 72768 VSS nch l=0.04u w=0.24u
m10168 5507 5510 5511 VSS nch l=0.13u w=1.3u
m10169 72781 5784 72765 VSS nch l=0.25u w=0.5u
m10170 72782 5732 72766 VSS nch l=0.25u w=0.5u
m10171 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10172 5749 4791 VSS VSS nch l=0.04u w=0.4u
m10173 5750 5746 VSS VSS nch l=0.04u w=0.4u
m10174 72785 5627 VSS VSS nch l=0.04u w=0.8u
m10175 72786 5748 VSS VSS nch l=0.04u w=0.8u
m10176 72788 5784 72774 VSS nch l=0.25u w=0.5u
m10177 72789 5784 72775 VSS nch l=0.25u w=0.5u
m10178 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10179 5751 5747 72785 VSS nch l=0.04u w=0.8u
m10180 5752 5869 72786 VSS nch l=0.04u w=0.8u
m10181 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10182 VSS 5784 72781 VSS nch l=0.25u w=0.5u
m10183 VSS 5732 72782 VSS nch l=0.25u w=0.5u
m10184 72797 4791 VSS VSS nch l=0.04u w=0.8u
m10185 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10186 5488 5784 72788 VSS nch l=0.25u w=0.5u
m10187 5488 5784 72789 VSS nch l=0.25u w=0.5u
m10188 72799 5750 VSS VSS nch l=0.04u w=0.8u
m10189 5765 4705 72797 VSS nch l=0.04u w=0.8u
m10190 5766 5525 5751 VSS nch l=0.04u w=0.4u
m10191 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10192 5767 5752 VSS VSS nch l=0.04u w=0.4u
m10193 5708 5797 72799 VSS nch l=0.04u w=0.8u
m10194 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10195 72810 5728 5766 VSS nch l=0.04u w=0.12u
m10196 VSS 5752 5767 VSS nch l=0.04u w=0.4u
m10197 72811 5784 5488 VSS nch l=0.25u w=0.5u
m10198 72812 5784 5488 VSS nch l=0.25u w=0.5u
m10199 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10200 VSS 5794 72810 VSS nch l=0.04u w=0.12u
m10201 72815 5749 VSS VSS nch l=0.04u w=0.8u
m10202 72821 5784 VSS VSS nch l=0.25u w=0.5u
m10203 72822 5784 VSS VSS nch l=0.25u w=0.5u
m10204 72823 5784 VSS VSS nch l=0.25u w=0.5u
m10205 72824 5784 VSS VSS nch l=0.25u w=0.5u
m10206 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10207 5770 5277 5750 VSS nch l=0.04u w=0.4u
m10208 72826 5784 72811 VSS nch l=0.25u w=0.5u
m10209 72827 5784 72812 VSS nch l=0.25u w=0.5u
m10210 5772 5766 VSS VSS nch l=0.04u w=0.4u
m10211 5768 5730 72815 VSS nch l=0.04u w=0.8u
m10212 5773 5836 VSS VSS nch l=0.04u w=0.4u
m10213 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10214 72828 5257 5770 VSS nch l=0.04u w=0.12u
m10215 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10216 72830 5784 72821 VSS nch l=0.25u w=0.5u
m10217 72831 5784 72822 VSS nch l=0.25u w=0.5u
m10218 5784 5814 5769 VSS nch l=0.25u w=0.65u
m10219 72832 5784 72823 VSS nch l=0.25u w=0.5u
m10220 72833 5784 72824 VSS nch l=0.25u w=0.5u
m10221 VSS 5790 72828 VSS nch l=0.04u w=0.12u
m10222 72834 5784 72826 VSS nch l=0.25u w=0.5u
m10223 72835 5784 72827 VSS nch l=0.25u w=0.5u
m10224 5339 5015 VDDREF VSS nch l=0.04u w=1.3u
m10225 72836 5627 VSS VSS nch l=0.04u w=0.8u
m10226 72838 5768 VSS VSS nch l=0.04u w=0.8u
m10227 VSS POSTDIV1[0] 5785 VSS nch l=0.04u w=0.8u
m10228 5790 5770 VSS VSS nch l=0.04u w=0.4u
m10229 VDDREF 5015 5339 VSS nch l=0.04u w=1.3u
m10230 5787 5772 72836 VSS nch l=0.04u w=0.8u
m10231 5769 5814 5784 VSS nch l=0.25u w=0.65u
m10232 5788 5765 72838 VSS nch l=0.04u w=0.8u
m10233 72842 5784 72830 VSS nch l=0.25u w=0.5u
m10234 72843 5784 72831 VSS nch l=0.25u w=0.5u
m10235 72844 5784 72832 VSS nch l=0.25u w=0.5u
m10236 72845 5784 72833 VSS nch l=0.25u w=0.5u
m10237 5785 POSTDIV1[0] VSS VSS nch l=0.04u w=0.8u
m10238 VSS 5784 72834 VSS nch l=0.25u w=0.5u
m10239 VSS 5784 72835 VSS nch l=0.25u w=0.5u
m10240 72850 5765 5788 VSS nch l=0.04u w=0.8u
m10241 5789 5773 5785 VSS nch l=0.04u w=0.62u
m10242 5793 5257 5790 VSS nch l=0.04u w=0.4u
m10243 5792 5784 72842 VSS nch l=0.25u w=0.5u
m10244 5792 5784 72843 VSS nch l=0.25u w=0.5u
m10245 5769 5784 72844 VSS nch l=0.25u w=0.5u
m10246 5769 5784 72845 VSS nch l=0.25u w=0.5u
m10247 VSS 5768 72850 VSS nch l=0.04u w=0.8u
m10248 5794 5787 VSS VSS nch l=0.04u w=0.4u
m10249 72857 5784 VSS VSS nch l=0.25u w=0.5u
m10250 72858 5784 VSS VSS nch l=0.25u w=0.5u
m10251 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10252 72859 5277 5793 VSS nch l=0.04u w=0.12u
m10253 72866 5789 VSS VSS nch l=0.04u w=0.8u
m10254 72867 5784 5769 VSS nch l=0.25u w=0.5u
m10255 72868 5784 5769 VSS nch l=0.25u w=0.5u
m10256 VSS 5797 72859 VSS nch l=0.04u w=0.12u
m10257 5796 BYPASS VSS VSS nch l=0.04u w=0.4u
m10258 72877 5784 72857 VSS nch l=0.25u w=0.5u
m10259 72878 5784 72858 VSS nch l=0.25u w=0.5u
m10260 5795 5824 72866 VSS nch l=0.04u w=0.8u
m10261 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10262 5797 5793 VSS VSS nch l=0.04u w=0.4u
m10263 VSS 4953 5627 VSS nch l=0.04u w=0.4u
m10264 72884 5784 72867 VSS nch l=0.25u w=0.5u
m10265 72885 5784 72868 VSS nch l=0.25u w=0.5u
m10266 5784 5814 5769 VSS nch l=0.25u w=0.65u
m10267 72888 5784 72877 VSS nch l=0.25u w=0.5u
m10268 72889 5784 72878 VSS nch l=0.25u w=0.5u
m10269 72890 5796 VSS VSS nch l=0.04u w=0.8u
m10270 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10271 72895 5824 5798 VSS nch l=0.04u w=0.8u
m10272 5799 PD 72890 VSS nch l=0.04u w=0.8u
m10273 5801 5790 VSS VSS nch l=0.04u w=0.4u
m10274 5802 FOUT1PH0 VSS VSS nch l=0.04u w=0.4u
m10275 72904 5814 VSS VSS nch l=0.25u w=0.5u
m10276 5769 5814 5784 VSS nch l=0.25u w=0.65u
m10277 72905 5784 72884 VSS nch l=0.25u w=0.5u
m10278 72906 5784 72885 VSS nch l=0.25u w=0.5u
m10279 72907 5807 72895 VSS nch l=0.04u w=0.8u
m10280 5488 5784 72888 VSS nch l=0.25u w=0.5u
m10281 5488 5784 72889 VSS nch l=0.25u w=0.5u
m10282 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10283 VSS FOUT1PH0 5802 VSS nch l=0.04u w=0.4u
m10284 VSS 4933 72907 VSS nch l=0.04u w=0.8u
m10285 72917 5799 VSS VSS nch l=0.04u w=0.8u
m10286 72918 5797 VSS VSS nch l=0.04u w=0.8u
m10287 5802 FOUT1PH0 VSS VSS nch l=0.04u w=0.4u
m10288 72919 5814 72904 VSS nch l=0.25u w=0.5u
m10289 VSS 5784 72905 VSS nch l=0.25u w=0.5u
m10290 VSS 5784 72906 VSS nch l=0.25u w=0.5u
m10291 72920 5784 5488 VSS nch l=0.25u w=0.5u
m10292 72921 5784 5488 VSS nch l=0.25u w=0.5u
m10293 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10294 5805 4703 72917 VSS nch l=0.04u w=0.8u
m10295 5806 5801 72918 VSS nch l=0.04u w=0.8u
m10296 VSS FOUT1PH0 5802 VSS nch l=0.04u w=0.4u
m10297 5808 5831 5807 VSS nch l=0.04u w=0.62u
m10298 72934 5784 VSS VSS nch l=0.25u w=0.5u
m10299 72935 5784 VSS VSS nch l=0.25u w=0.5u
m10300 72936 5814 72919 VSS nch l=0.25u w=0.5u
m10301 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10302 72937 5784 72920 VSS nch l=0.25u w=0.5u
m10303 72938 5784 72921 VSS nch l=0.25u w=0.5u
m10304 VSS POSTDIV1[0] 5808 VSS nch l=0.04u w=0.8u
m10305 VSS 5788 5811 VSS nch l=0.04u w=0.4u
m10306 VSS 5806 5812 VSS nch l=0.04u w=0.4u
m10307 VSS 5363 5813 VSS nch l=0.04u w=0.4u
m10308 5808 POSTDIV1[0] VSS VSS nch l=0.04u w=0.8u
m10309 5783 5814 5810 VSS nch l=0.25u w=0.65u
m10310 72947 5784 72934 VSS nch l=0.25u w=0.5u
m10311 72948 5784 72935 VSS nch l=0.25u w=0.5u
m10312 5814 5814 72936 VSS nch l=0.25u w=0.5u
m10313 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10314 5817 5811 VSS VSS nch l=0.04u w=0.4u
m10315 5818 5812 VSS VSS nch l=0.04u w=0.4u
m10316 5819 5813 VSS VSS nch l=0.04u w=0.4u
m10317 72953 5784 72937 VSS nch l=0.25u w=0.5u
m10318 72954 5784 72938 VSS nch l=0.25u w=0.5u
m10319 5810 5814 5783 VSS nch l=0.25u w=0.65u
m10320 72960 5784 72947 VSS nch l=0.25u w=0.5u
m10321 72961 5784 72948 VSS nch l=0.25u w=0.5u
m10322 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10323 VSS 5784 72953 VSS nch l=0.25u w=0.5u
m10324 VSS 5784 72954 VSS nch l=0.25u w=0.5u
m10325 VSS 5901 5820 VSS nch l=0.04u w=0.8u
m10326 VSS 5902 5821 VSS nch l=0.04u w=0.8u
m10327 VSS 5903 5822 VSS nch l=0.04u w=0.8u
m10328 VSS 5829 5824 VSS nch l=0.04u w=0.4u
m10329 5820 5901 VSS VSS nch l=0.04u w=0.8u
m10330 5821 5902 VSS VSS nch l=0.04u w=0.8u
m10331 5822 5903 VSS VSS nch l=0.04u w=0.8u
m10332 72973 5824 VSS VSS nch l=0.04u w=0.12u
m10333 5810 5784 72960 VSS nch l=0.25u w=0.5u
m10334 5810 5784 72961 VSS nch l=0.25u w=0.5u
m10335 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10336 5825 5788 5820 VSS nch l=0.04u w=0.8u
m10337 5826 5806 5821 VSS nch l=0.04u w=0.8u
m10338 5827 5363 5822 VSS nch l=0.04u w=0.8u
m10339 5829 5837 72973 VSS nch l=0.04u w=0.12u
m10340 72981 5784 5810 VSS nch l=0.25u w=0.5u
m10341 72982 5784 5810 VSS nch l=0.25u w=0.5u
m10342 5339 5814 5488 VSS nch l=0.25u w=0.65u
m10343 5339 5814 5488 VSS nch l=0.25u w=0.65u
m10344 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10345 72983 5784 5792 VSS nch l=0.25u w=0.5u
m10346 72984 5784 5792 VSS nch l=0.25u w=0.5u
m10347 5831 5864 5829 VSS nch l=0.04u w=0.4u
m10348 FOUTPOSTDIV 5825 VSS VSS nch l=0.04u w=0.4u
m10349 FOUT3 5826 VSS VSS nch l=0.04u w=0.4u
m10350 FOUT1PH0 5827 VSS VSS nch l=0.04u w=0.4u
m10351 5488 5814 5339 VSS nch l=0.25u w=0.65u
m10352 5488 5814 5339 VSS nch l=0.25u w=0.65u
m10353 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10354 72989 5784 72981 VSS nch l=0.25u w=0.5u
m10355 72990 5784 72982 VSS nch l=0.25u w=0.5u
m10356 VSS 5825 FOUTPOSTDIV VSS nch l=0.04u w=0.4u
m10357 VSS 5826 FOUT3 VSS nch l=0.04u w=0.4u
m10358 VSS 5827 FOUT1PH0 VSS nch l=0.04u w=0.4u
m10359 72992 5784 72983 VSS nch l=0.25u w=0.5u
m10360 72993 5784 72984 VSS nch l=0.25u w=0.5u
m10361 5783 5814 5810 VSS nch l=0.25u w=0.65u
m10362 VSS 5835 5831 VSS nch l=0.04u w=0.4u
m10363 FOUTPOSTDIV 5825 VSS VSS nch l=0.04u w=0.4u
m10364 FOUT3 5826 VSS VSS nch l=0.04u w=0.4u
m10365 FOUT1PH0 5827 VSS VSS nch l=0.04u w=0.4u
m10366 72999 5831 VSS VSS nch l=0.04u w=0.12u
m10367 5339 5814 5488 VSS nch l=0.25u w=0.65u
m10368 5339 5814 5488 VSS nch l=0.25u w=0.65u
m10369 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10370 5810 5814 5783 VSS nch l=0.25u w=0.65u
m10371 73000 5784 72989 VSS nch l=0.25u w=0.5u
m10372 73001 5784 72990 VSS nch l=0.25u w=0.5u
m10373 73002 5784 72992 VSS nch l=0.25u w=0.5u
m10374 73003 5784 72993 VSS nch l=0.25u w=0.5u
m10375 VSS 5825 FOUTPOSTDIV VSS nch l=0.04u w=0.4u
m10376 VSS 5826 FOUT3 VSS nch l=0.04u w=0.4u
m10377 VSS 5827 FOUT1PH0 VSS nch l=0.04u w=0.4u
m10378 5835 5864 72999 VSS nch l=0.04u w=0.12u
m10379 FOUTPOSTDIV 5825 VSS VSS nch l=0.04u w=0.4u
m10380 FOUT3 5826 VSS VSS nch l=0.04u w=0.4u
m10381 FOUT1PH0 5827 VSS VSS nch l=0.04u w=0.4u
m10382 5488 5814 5339 VSS nch l=0.25u w=0.65u
m10383 5488 5814 5339 VSS nch l=0.25u w=0.65u
m10384 VSS 5015 VSS VSS nch l=0.25u w=1.3u
m10385 5836 5837 5835 VSS nch l=0.04u w=0.4u
m10386 VSS 5784 73000 VSS nch l=0.25u w=0.5u
m10387 VSS 5784 73001 VSS nch l=0.25u w=0.5u
m10388 VSS 5784 73002 VSS nch l=0.25u w=0.5u
m10389 VSS 5784 73003 VSS nch l=0.25u w=0.5u
m10390 VSS 5825 FOUTPOSTDIV VSS nch l=0.04u w=0.4u
m10391 VSS 5826 FOUT3 VSS nch l=0.04u w=0.4u
m10392 VSS 5827 FOUT1PH0 VSS nch l=0.04u w=0.4u
m10393 FOUTPOSTDIV 5825 VSS VSS nch l=0.04u w=0.4u
m10394 FOUT3 5826 VSS VSS nch l=0.04u w=0.4u
m10395 FOUT1PH0 5827 VSS VSS nch l=0.04u w=0.4u
m10396 VSS 5864 5837 VSS nch l=0.04u w=0.4u
m10397 VSS 5825 FOUTPOSTDIV VSS nch l=0.04u w=0.4u
m10398 VSS 5826 FOUT3 VSS nch l=0.04u w=0.4u
m10399 VSS 5827 FOUT1PH0 VSS nch l=0.04u w=0.4u
m10400 VSS 5844 5836 VSS nch l=0.04u w=0.4u
m10401 VSS 5817 5838 VSS nch l=0.04u w=0.4u
m10402 VSS 5818 5839 VSS nch l=0.04u w=0.4u
m10403 VSS 5819 5840 VSS nch l=0.04u w=0.4u
m10404 73038 5836 VSS VSS nch l=0.04u w=0.12u
m10405 5844 5859 73038 VSS nch l=0.04u w=0.12u
m10406 5845 5838 5841 VSS nch l=0.04u w=0.4u
m10407 5846 5839 5842 VSS nch l=0.04u w=0.4u
m10408 5847 5840 5843 VSS nch l=0.04u w=0.4u
m10409 5848 5864 5844 VSS nch l=0.04u w=0.4u
m10410 73044 5817 5845 VSS nch l=0.04u w=0.24u
m10411 73045 5818 5846 VSS nch l=0.04u w=0.24u
m10412 73046 5819 5847 VSS nch l=0.04u w=0.24u
m10413 VSS 5849 73044 VSS nch l=0.04u w=0.24u
m10414 VSS 5850 73045 VSS nch l=0.04u w=0.24u
m10415 VSS 5851 73046 VSS nch l=0.04u w=0.24u
m10416 VSS 5853 5848 VSS nch l=0.04u w=0.4u
m10417 73051 5841 VSS VSS nch l=0.04u w=0.8u
m10418 73052 5842 VSS VSS nch l=0.04u w=0.8u
m10419 73053 5843 VSS VSS nch l=0.04u w=0.8u
m10420 73055 5848 VSS VSS nch l=0.04u w=0.12u
m10421 5849 5845 73051 VSS nch l=0.04u w=0.8u
m10422 5850 5846 73052 VSS nch l=0.04u w=0.8u
m10423 5851 5847 73053 VSS nch l=0.04u w=0.8u
m10424 5853 5864 73055 VSS nch l=0.04u w=0.12u
m10425 5795 5859 5853 VSS nch l=0.04u w=0.4u
m10426 5855 5817 5849 VSS nch l=0.04u w=0.4u
m10427 5856 5818 5850 VSS nch l=0.04u w=0.4u
m10428 5857 5819 5851 VSS nch l=0.04u w=0.4u
m10429 73118 5838 5855 VSS nch l=0.04u w=0.12u
m10430 73119 5839 5856 VSS nch l=0.04u w=0.12u
m10431 73120 5840 5857 VSS nch l=0.04u w=0.12u
m10432 VSS 5864 5859 VSS nch l=0.04u w=0.4u
m10433 VSS 5870 73118 VSS nch l=0.04u w=0.12u
m10434 VSS 5871 73119 VSS nch l=0.04u w=0.12u
m10435 VSS 5872 73120 VSS nch l=0.04u w=0.12u
m10436 5861 5855 VSS VSS nch l=0.04u w=0.4u
m10437 5862 5856 VSS VSS nch l=0.04u w=0.4u
m10438 5863 5857 VSS VSS nch l=0.04u w=0.4u
m10439 5865 4708 5864 VSS nch l=0.04u w=0.8u
m10440 73140 5841 VSS VSS nch l=0.04u w=0.8u
m10441 73141 5842 VSS VSS nch l=0.04u w=0.8u
m10442 73142 5843 VSS VSS nch l=0.04u w=0.8u
m10443 VSS 4933 5865 VSS nch l=0.04u w=0.8u
m10444 5866 5861 73140 VSS nch l=0.04u w=0.8u
m10445 5867 5862 73141 VSS nch l=0.04u w=0.8u
m10446 5868 5863 73142 VSS nch l=0.04u w=0.8u
m10447 5865 4933 VSS VSS nch l=0.04u w=0.8u
m10448 5870 5866 VSS VSS nch l=0.04u w=0.4u
m10449 5871 5867 VSS VSS nch l=0.04u w=0.4u
m10450 5872 5868 VSS VSS nch l=0.04u w=0.4u
m10451 5873 5877 5869 VSS nch l=0.04u w=0.62u
m10452 VSS 4925 5873 VSS nch l=0.04u w=0.8u
m10453 VSS 5817 5874 VSS nch l=0.04u w=0.4u
m10454 VSS 5818 5875 VSS nch l=0.04u w=0.4u
m10455 VSS 5819 5876 VSS nch l=0.04u w=0.4u
m10456 5873 4925 VSS VSS nch l=0.04u w=0.8u
m10457 5878 5874 5870 VSS nch l=0.04u w=0.4u
m10458 5879 5875 5871 VSS nch l=0.04u w=0.4u
m10459 5880 5876 5872 VSS nch l=0.04u w=0.4u
m10460 VSS 5881 5877 VSS nch l=0.04u w=0.4u
m10461 73184 5817 5878 VSS nch l=0.04u w=0.24u
m10462 73185 5818 5879 VSS nch l=0.04u w=0.24u
m10463 73186 5819 5880 VSS nch l=0.04u w=0.24u
m10464 73188 5877 VSS VSS nch l=0.04u w=0.12u
m10465 VSS 5883 73184 VSS nch l=0.04u w=0.24u
m10466 VSS 5884 73185 VSS nch l=0.04u w=0.24u
m10467 VSS 5885 73186 VSS nch l=0.04u w=0.24u
m10468 5881 5895 73188 VSS nch l=0.04u w=0.12u
m10469 73192 5841 VSS VSS nch l=0.04u w=0.8u
m10470 73193 5842 VSS VSS nch l=0.04u w=0.8u
m10471 73194 5843 VSS VSS nch l=0.04u w=0.8u
m10472 5886 5899 5881 VSS nch l=0.04u w=0.4u
m10473 5883 5878 73192 VSS nch l=0.04u w=0.8u
m10474 5884 5879 73193 VSS nch l=0.04u w=0.8u
m10475 5885 5880 73194 VSS nch l=0.04u w=0.8u
m10476 VSS 5890 5886 VSS nch l=0.04u w=0.4u
m10477 5887 5817 5883 VSS nch l=0.04u w=0.4u
m10478 5888 5818 5884 VSS nch l=0.04u w=0.4u
m10479 5889 5819 5885 VSS nch l=0.04u w=0.4u
m10480 73198 5886 VSS VSS nch l=0.04u w=0.12u
m10481 73199 5874 5887 VSS nch l=0.04u w=0.12u
m10482 73200 5875 5888 VSS nch l=0.04u w=0.12u
m10483 73201 5876 5889 VSS nch l=0.04u w=0.12u
m10484 5890 5899 73198 VSS nch l=0.04u w=0.12u
m10485 VSS 5901 73199 VSS nch l=0.04u w=0.12u
m10486 VSS 5902 73200 VSS nch l=0.04u w=0.12u
m10487 VSS 5903 73201 VSS nch l=0.04u w=0.12u
m10488 5891 5895 5890 VSS nch l=0.04u w=0.4u
m10489 5892 5887 VSS VSS nch l=0.04u w=0.4u
m10490 5893 5888 VSS VSS nch l=0.04u w=0.4u
m10491 5894 5889 VSS VSS nch l=0.04u w=0.4u
m10492 VSS 5899 5895 VSS nch l=0.04u w=0.4u
m10493 73202 5841 VSS VSS nch l=0.04u w=0.8u
m10494 73203 5842 VSS VSS nch l=0.04u w=0.8u
m10495 73204 5843 VSS VSS nch l=0.04u w=0.8u
m10496 5896 5892 73202 VSS nch l=0.04u w=0.8u
m10497 5897 5893 73203 VSS nch l=0.04u w=0.8u
m10498 5898 5894 73204 VSS nch l=0.04u w=0.8u
m10499 5900 4708 5899 VSS nch l=0.04u w=0.62u
m10500 5901 5896 VSS VSS nch l=0.04u w=0.4u
m10501 5902 5897 VSS VSS nch l=0.04u w=0.4u
m10502 5903 5898 VSS VSS nch l=0.04u w=0.4u
m10503 VSS 4925 5900 VSS nch l=0.04u w=0.8u
m10504 5900 4925 VSS VSS nch l=0.04u w=0.8u
m10505 VSS 5877 5891 VSS nch l=0.04u w=0.4u
m10506 VSS 5805 5841 VSS nch l=0.04u w=0.4u
m10507 VSS 4953 5842 VSS nch l=0.04u w=0.4u
m10508 VSS 4953 5843 VSS nch l=0.04u w=0.4u
m10509 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10510 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10511 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10512 4737 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10513 4738 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10514 4749 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10515 4750 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10516 4761 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10517 4762 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10518 4773 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10519 4774 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10520 4785 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10521 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10522 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10523 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10524 4737 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10525 4738 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10526 4749 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10527 4750 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10528 4761 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10529 4762 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10530 4773 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10531 4774 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10532 4785 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10533 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10534 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10535 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10536 4737 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10537 4738 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10538 4749 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10539 4750 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10540 4761 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10541 4762 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10542 4773 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10543 4774 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10544 4785 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10545 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10546 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10547 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10548 4737 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10549 4738 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10550 4749 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10551 4750 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10552 4761 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10553 4762 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10554 4773 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10555 4774 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10556 4785 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10557 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10558 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10559 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10560 4737 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10561 4738 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10562 4749 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10563 4750 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10564 4761 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10565 4762 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10566 4773 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10567 4774 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10568 4785 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10569 4797 5643 5002 VDDHV pch_18 l=0.27u w=1.66u
m10570 4806 5643 5003 VDDHV pch_18 l=0.27u w=1.66u
m10571 4807 5643 5004 VDDHV pch_18 l=0.27u w=1.66u
m10572 4816 5643 5005 VDDHV pch_18 l=0.27u w=1.66u
m10573 4817 5643 5006 VDDHV pch_18 l=0.27u w=1.66u
m10574 4826 5643 5007 VDDHV pch_18 l=0.27u w=1.66u
m10575 4827 5643 5008 VDDHV pch_18 l=0.27u w=1.66u
m10576 4836 5643 5009 VDDHV pch_18 l=0.27u w=1.66u
m10577 4837 5643 5010 VDDHV pch_18 l=0.27u w=1.66u
m10578 4846 5643 5011 VDDHV pch_18 l=0.27u w=1.66u
m10579 4847 5643 5012 VDDHV pch_18 l=0.27u w=1.66u
m10580 4856 5643 5013 VDDHV pch_18 l=0.27u w=1.66u
m10581 4717 5643 5025 VDDHV pch_18 l=0.27u w=1.66u
m10582 4726 5643 5026 VDDHV pch_18 l=0.27u w=1.66u
m10583 4727 5643 5027 VDDHV pch_18 l=0.27u w=1.66u
m10584 4736 5643 5028 VDDHV pch_18 l=0.27u w=1.66u
m10585 4739 5643 5029 VDDHV pch_18 l=0.27u w=1.66u
m10586 4748 5643 5030 VDDHV pch_18 l=0.27u w=1.66u
m10587 4751 5643 5031 VDDHV pch_18 l=0.27u w=1.66u
m10588 4760 5643 5032 VDDHV pch_18 l=0.27u w=1.66u
m10589 4763 5643 5033 VDDHV pch_18 l=0.27u w=1.66u
m10590 4772 5643 5034 VDDHV pch_18 l=0.27u w=1.66u
m10591 4775 5643 5035 VDDHV pch_18 l=0.27u w=1.66u
m10592 4784 5643 5036 VDDHV pch_18 l=0.27u w=1.66u
m10593 4718 5643 5052 VDDHV pch_18 l=0.27u w=1.66u
m10594 4725 5643 5053 VDDHV pch_18 l=0.27u w=1.66u
m10595 4728 5643 5054 VDDHV pch_18 l=0.27u w=1.66u
m10596 4735 5643 5055 VDDHV pch_18 l=0.27u w=1.66u
m10597 4740 5643 5056 VDDHV pch_18 l=0.27u w=1.66u
m10598 4747 5643 5057 VDDHV pch_18 l=0.27u w=1.66u
m10599 4752 5643 5058 VDDHV pch_18 l=0.27u w=1.66u
m10600 4759 5643 5059 VDDHV pch_18 l=0.27u w=1.66u
m10601 4764 5643 5060 VDDHV pch_18 l=0.27u w=1.66u
m10602 4771 5643 5061 VDDHV pch_18 l=0.27u w=1.66u
m10603 4776 5643 5062 VDDHV pch_18 l=0.27u w=1.66u
m10604 4783 5643 5063 VDDHV pch_18 l=0.27u w=1.66u
m10605 4798 5643 5073 VDDHV pch_18 l=0.27u w=1.66u
m10606 4805 5643 5074 VDDHV pch_18 l=0.27u w=1.66u
m10607 4808 5643 5075 VDDHV pch_18 l=0.27u w=1.66u
m10608 4815 5643 5076 VDDHV pch_18 l=0.27u w=1.66u
m10609 4818 5643 5077 VDDHV pch_18 l=0.27u w=1.66u
m10610 4825 5643 5078 VDDHV pch_18 l=0.27u w=1.66u
m10611 4828 5643 5079 VDDHV pch_18 l=0.27u w=1.66u
m10612 4835 5643 5080 VDDHV pch_18 l=0.27u w=1.66u
m10613 4838 5643 5081 VDDHV pch_18 l=0.27u w=1.66u
m10614 4845 5643 5082 VDDHV pch_18 l=0.27u w=1.66u
m10615 4848 5643 5083 VDDHV pch_18 l=0.27u w=1.66u
m10616 4855 5643 5084 VDDHV pch_18 l=0.27u w=1.66u
m10617 4877 5643 5098 VDDHV pch_18 l=0.27u w=1.66u
m10618 4884 5643 5099 VDDHV pch_18 l=0.27u w=1.66u
m10619 4885 5643 5100 VDDHV pch_18 l=0.27u w=1.66u
m10620 4892 5643 5101 VDDHV pch_18 l=0.27u w=1.66u
m10621 4893 5643 5102 VDDHV pch_18 l=0.27u w=1.66u
m10622 4900 5643 5103 VDDHV pch_18 l=0.27u w=1.66u
m10623 4901 5643 5104 VDDHV pch_18 l=0.27u w=1.66u
m10624 4908 5643 5105 VDDHV pch_18 l=0.27u w=1.66u
m10625 4909 5643 5106 VDDHV pch_18 l=0.27u w=1.66u
m10626 4916 5643 5107 VDDHV pch_18 l=0.27u w=1.66u
m10627 4917 5643 5108 VDDHV pch_18 l=0.27u w=1.66u
m10628 4924 5643 5109 VDDHV pch_18 l=0.27u w=1.66u
m10629 4878 5643 5118 VDDHV pch_18 l=0.27u w=1.66u
m10630 4883 5643 5119 VDDHV pch_18 l=0.27u w=1.66u
m10631 4886 5643 5120 VDDHV pch_18 l=0.27u w=1.66u
m10632 4891 5643 5121 VDDHV pch_18 l=0.27u w=1.66u
m10633 4894 5643 5122 VDDHV pch_18 l=0.27u w=1.66u
m10634 4899 5643 5123 VDDHV pch_18 l=0.27u w=1.66u
m10635 4902 5643 5124 VDDHV pch_18 l=0.27u w=1.66u
m10636 4907 5643 5125 VDDHV pch_18 l=0.27u w=1.66u
m10637 4910 5643 5126 VDDHV pch_18 l=0.27u w=1.66u
m10638 4915 5643 5127 VDDHV pch_18 l=0.27u w=1.66u
m10639 4918 5643 5128 VDDHV pch_18 l=0.27u w=1.66u
m10640 4923 5643 5129 VDDHV pch_18 l=0.27u w=1.66u
m10641 4799 5643 5144 VDDHV pch_18 l=0.27u w=1.66u
m10642 4804 5643 5145 VDDHV pch_18 l=0.27u w=1.66u
m10643 4809 5643 5146 VDDHV pch_18 l=0.27u w=1.66u
m10644 4814 5643 5147 VDDHV pch_18 l=0.27u w=1.66u
m10645 4819 5643 5148 VDDHV pch_18 l=0.27u w=1.66u
m10646 4824 5643 5149 VDDHV pch_18 l=0.27u w=1.66u
m10647 4829 5643 5150 VDDHV pch_18 l=0.27u w=1.66u
m10648 4834 5643 5151 VDDHV pch_18 l=0.27u w=1.66u
m10649 4839 5643 5152 VDDHV pch_18 l=0.27u w=1.66u
m10650 4844 5643 5153 VDDHV pch_18 l=0.27u w=1.66u
m10651 4849 5643 5154 VDDHV pch_18 l=0.27u w=1.66u
m10652 4854 5643 5155 VDDHV pch_18 l=0.27u w=1.66u
m10653 4719 5643 5165 VDDHV pch_18 l=0.27u w=1.66u
m10654 4724 5643 5166 VDDHV pch_18 l=0.27u w=1.66u
m10655 4729 5643 5167 VDDHV pch_18 l=0.27u w=1.66u
m10656 4734 5643 5168 VDDHV pch_18 l=0.27u w=1.66u
m10657 4741 5643 5169 VDDHV pch_18 l=0.27u w=1.66u
m10658 4746 5643 5170 VDDHV pch_18 l=0.27u w=1.66u
m10659 4753 5643 5171 VDDHV pch_18 l=0.27u w=1.66u
m10660 4758 5643 5172 VDDHV pch_18 l=0.27u w=1.66u
m10661 4765 5643 5173 VDDHV pch_18 l=0.27u w=1.66u
m10662 4770 5643 5174 VDDHV pch_18 l=0.27u w=1.66u
m10663 4777 5643 5175 VDDHV pch_18 l=0.27u w=1.66u
m10664 4782 5643 5176 VDDHV pch_18 l=0.27u w=1.66u
m10665 4720 5643 5191 VDDHV pch_18 l=0.27u w=1.66u
m10666 4723 5643 5192 VDDHV pch_18 l=0.27u w=1.66u
m10667 4730 5643 5193 VDDHV pch_18 l=0.27u w=1.66u
m10668 4733 5643 5194 VDDHV pch_18 l=0.27u w=1.66u
m10669 4742 5643 5195 VDDHV pch_18 l=0.27u w=1.66u
m10670 4745 5643 5196 VDDHV pch_18 l=0.27u w=1.66u
m10671 4754 5643 5197 VDDHV pch_18 l=0.27u w=1.66u
m10672 4757 5643 5198 VDDHV pch_18 l=0.27u w=1.66u
m10673 4766 5643 5199 VDDHV pch_18 l=0.27u w=1.66u
m10674 4769 5643 5200 VDDHV pch_18 l=0.27u w=1.66u
m10675 4778 5643 5201 VDDHV pch_18 l=0.27u w=1.66u
m10676 4781 5643 5202 VDDHV pch_18 l=0.27u w=1.66u
m10677 4800 5643 5214 VDDHV pch_18 l=0.27u w=1.66u
m10678 4803 5643 5215 VDDHV pch_18 l=0.27u w=1.66u
m10679 4810 5643 5216 VDDHV pch_18 l=0.27u w=1.66u
m10680 4813 5643 5217 VDDHV pch_18 l=0.27u w=1.66u
m10681 4820 5643 5218 VDDHV pch_18 l=0.27u w=1.66u
m10682 4823 5643 5219 VDDHV pch_18 l=0.27u w=1.66u
m10683 4830 5643 5220 VDDHV pch_18 l=0.27u w=1.66u
m10684 4833 5643 5221 VDDHV pch_18 l=0.27u w=1.66u
m10685 4840 5643 5222 VDDHV pch_18 l=0.27u w=1.66u
m10686 4843 5643 5223 VDDHV pch_18 l=0.27u w=1.66u
m10687 4850 5643 5224 VDDHV pch_18 l=0.27u w=1.66u
m10688 4853 5643 5225 VDDHV pch_18 l=0.27u w=1.66u
m10689 4879 5643 5236 VDDHV pch_18 l=0.27u w=1.66u
m10690 4882 5643 5237 VDDHV pch_18 l=0.27u w=1.66u
m10691 4887 5643 5238 VDDHV pch_18 l=0.27u w=1.66u
m10692 4890 5643 5239 VDDHV pch_18 l=0.27u w=1.66u
m10693 4895 5643 5240 VDDHV pch_18 l=0.27u w=1.66u
m10694 4898 5643 5241 VDDHV pch_18 l=0.27u w=1.66u
m10695 4903 5643 5242 VDDHV pch_18 l=0.27u w=1.66u
m10696 4906 5643 5243 VDDHV pch_18 l=0.27u w=1.66u
m10697 4911 5643 5244 VDDHV pch_18 l=0.27u w=1.66u
m10698 4914 5643 5245 VDDHV pch_18 l=0.27u w=1.66u
m10699 4919 5643 5246 VDDHV pch_18 l=0.27u w=1.66u
m10700 4922 5643 5247 VDDHV pch_18 l=0.27u w=1.66u
m10701 4880 5643 5258 VDDHV pch_18 l=0.27u w=1.66u
m10702 4881 5643 5259 VDDHV pch_18 l=0.27u w=1.66u
m10703 4888 5643 5260 VDDHV pch_18 l=0.27u w=1.66u
m10704 4889 5643 5261 VDDHV pch_18 l=0.27u w=1.66u
m10705 4896 5643 5262 VDDHV pch_18 l=0.27u w=1.66u
m10706 4897 5643 5263 VDDHV pch_18 l=0.27u w=1.66u
m10707 4904 5643 5264 VDDHV pch_18 l=0.27u w=1.66u
m10708 4905 5643 5265 VDDHV pch_18 l=0.27u w=1.66u
m10709 4912 5643 5266 VDDHV pch_18 l=0.27u w=1.66u
m10710 4913 5643 5267 VDDHV pch_18 l=0.27u w=1.66u
m10711 4920 5643 5268 VDDHV pch_18 l=0.27u w=1.66u
m10712 4921 5643 5269 VDDHV pch_18 l=0.27u w=1.66u
m10713 4801 5643 5279 VDDHV pch_18 l=0.27u w=1.66u
m10714 4802 5643 5280 VDDHV pch_18 l=0.27u w=1.66u
m10715 4811 5643 5281 VDDHV pch_18 l=0.27u w=1.66u
m10716 4812 5643 5282 VDDHV pch_18 l=0.27u w=1.66u
m10717 4821 5643 5283 VDDHV pch_18 l=0.27u w=1.66u
m10718 4822 5643 5284 VDDHV pch_18 l=0.27u w=1.66u
m10719 4831 5643 5285 VDDHV pch_18 l=0.27u w=1.66u
m10720 4832 5643 5286 VDDHV pch_18 l=0.27u w=1.66u
m10721 4841 5643 5287 VDDHV pch_18 l=0.27u w=1.66u
m10722 4842 5643 5288 VDDHV pch_18 l=0.27u w=1.66u
m10723 4851 5643 5289 VDDHV pch_18 l=0.27u w=1.66u
m10724 4852 5643 5290 VDDHV pch_18 l=0.27u w=1.66u
m10725 4721 5643 5298 VDDHV pch_18 l=0.27u w=1.66u
m10726 4722 5643 5299 VDDHV pch_18 l=0.27u w=1.66u
m10727 4731 5643 5300 VDDHV pch_18 l=0.27u w=1.66u
m10728 4732 5643 5301 VDDHV pch_18 l=0.27u w=1.66u
m10729 4743 5643 5302 VDDHV pch_18 l=0.27u w=1.66u
m10730 4744 5643 5303 VDDHV pch_18 l=0.27u w=1.66u
m10731 4755 5643 5304 VDDHV pch_18 l=0.27u w=1.66u
m10732 4756 5643 5305 VDDHV pch_18 l=0.27u w=1.66u
m10733 4767 5643 5306 VDDHV pch_18 l=0.27u w=1.66u
m10734 4768 5643 5307 VDDHV pch_18 l=0.27u w=1.66u
m10735 4779 5643 5308 VDDHV pch_18 l=0.27u w=1.66u
m10736 4780 5643 5309 VDDHV pch_18 l=0.27u w=1.66u
m10737 5344 5643 5325 VDDHV pch_18 l=0.27u w=1.66u
m10738 5345 5643 5326 VDDHV pch_18 l=0.27u w=1.66u
m10739 5346 5643 5327 VDDHV pch_18 l=0.27u w=1.66u
m10740 5347 5643 5328 VDDHV pch_18 l=0.27u w=1.66u
m10741 5348 5643 5329 VDDHV pch_18 l=0.27u w=1.66u
m10742 5349 5643 5330 VDDHV pch_18 l=0.27u w=1.66u
m10743 5350 5643 5331 VDDHV pch_18 l=0.27u w=1.66u
m10744 5351 5643 5332 VDDHV pch_18 l=0.27u w=1.66u
m10745 5352 5643 5333 VDDHV pch_18 l=0.27u w=1.66u
m10746 5353 5643 5334 VDDHV pch_18 l=0.27u w=1.66u
m10747 5354 5643 5335 VDDHV pch_18 l=0.27u w=1.66u
m10748 5355 5643 5336 VDDHV pch_18 l=0.27u w=1.66u
m10749 5380 5643 5365 VDDHV pch_18 l=0.27u w=1.66u
m10750 5381 5643 5366 VDDHV pch_18 l=0.27u w=1.66u
m10751 5382 5643 5367 VDDHV pch_18 l=0.27u w=1.66u
m10752 5383 5643 5368 VDDHV pch_18 l=0.27u w=1.66u
m10753 5384 5643 5369 VDDHV pch_18 l=0.27u w=1.66u
m10754 5385 5643 5370 VDDHV pch_18 l=0.27u w=1.66u
m10755 5386 5643 5371 VDDHV pch_18 l=0.27u w=1.66u
m10756 5387 5643 5372 VDDHV pch_18 l=0.27u w=1.66u
m10757 5388 5643 5373 VDDHV pch_18 l=0.27u w=1.66u
m10758 5389 5643 5374 VDDHV pch_18 l=0.27u w=1.66u
m10759 5390 5643 5375 VDDHV pch_18 l=0.27u w=1.66u
m10760 5391 5643 5376 VDDHV pch_18 l=0.27u w=1.66u
m10761 5411 5643 5397 VDDHV pch_18 l=0.27u w=1.66u
m10762 5412 5643 5398 VDDHV pch_18 l=0.27u w=1.66u
m10763 5413 5643 5399 VDDHV pch_18 l=0.27u w=1.66u
m10764 5414 5643 5400 VDDHV pch_18 l=0.27u w=1.66u
m10765 5415 5643 5401 VDDHV pch_18 l=0.27u w=1.66u
m10766 5416 5643 5402 VDDHV pch_18 l=0.27u w=1.66u
m10767 5417 5643 5403 VDDHV pch_18 l=0.27u w=1.66u
m10768 5418 5643 5404 VDDHV pch_18 l=0.27u w=1.66u
m10769 5419 5643 5405 VDDHV pch_18 l=0.27u w=1.66u
m10770 5420 5643 5406 VDDHV pch_18 l=0.27u w=1.66u
m10771 5421 5643 5407 VDDHV pch_18 l=0.27u w=1.66u
m10772 5422 5643 5408 VDDHV pch_18 l=0.27u w=1.66u
m10773 5442 5643 5427 VDDHV pch_18 l=0.27u w=1.66u
m10774 5443 5643 5428 VDDHV pch_18 l=0.27u w=1.66u
m10775 5444 5643 5429 VDDHV pch_18 l=0.27u w=1.66u
m10776 5445 5643 5430 VDDHV pch_18 l=0.27u w=1.66u
m10777 5446 5643 5431 VDDHV pch_18 l=0.27u w=1.66u
m10778 5447 5643 5432 VDDHV pch_18 l=0.27u w=1.66u
m10779 5448 5643 5433 VDDHV pch_18 l=0.27u w=1.66u
m10780 5449 5643 5434 VDDHV pch_18 l=0.27u w=1.66u
m10781 5450 5643 5435 VDDHV pch_18 l=0.27u w=1.66u
m10782 5451 5643 5436 VDDHV pch_18 l=0.27u w=1.66u
m10783 5452 5643 5437 VDDHV pch_18 l=0.27u w=1.66u
m10784 5453 5643 5438 VDDHV pch_18 l=0.27u w=1.66u
m10785 5474 5643 5459 VDDHV pch_18 l=0.27u w=1.66u
m10786 5475 5643 5460 VDDHV pch_18 l=0.27u w=1.66u
m10787 5476 5643 5461 VDDHV pch_18 l=0.27u w=1.66u
m10788 5477 5643 5462 VDDHV pch_18 l=0.27u w=1.66u
m10789 5478 5643 5463 VDDHV pch_18 l=0.27u w=1.66u
m10790 5479 5643 5464 VDDHV pch_18 l=0.27u w=1.66u
m10791 5480 5643 5465 VDDHV pch_18 l=0.27u w=1.66u
m10792 5481 5643 5466 VDDHV pch_18 l=0.27u w=1.66u
m10793 5482 5643 5467 VDDHV pch_18 l=0.27u w=1.66u
m10794 5483 5643 5468 VDDHV pch_18 l=0.27u w=1.66u
m10795 5484 5643 5469 VDDHV pch_18 l=0.27u w=1.66u
m10796 5485 5643 5470 VDDHV pch_18 l=0.27u w=1.66u
m10797 5506 5314 2 VDDHV pch_18 l=0.28u w=0.44u
m10798 5513 5643 5491 VDDHV pch_18 l=0.27u w=1.66u
m10799 5514 5643 5492 VDDHV pch_18 l=0.27u w=1.66u
m10800 5515 5643 5493 VDDHV pch_18 l=0.27u w=1.66u
m10801 5516 5643 5494 VDDHV pch_18 l=0.27u w=1.66u
m10802 5517 5643 5495 VDDHV pch_18 l=0.27u w=1.66u
m10803 5518 5643 5496 VDDHV pch_18 l=0.27u w=1.66u
m10804 5519 5643 5497 VDDHV pch_18 l=0.27u w=1.66u
m10805 5520 5643 5498 VDDHV pch_18 l=0.27u w=1.66u
m10806 5521 5643 5499 VDDHV pch_18 l=0.27u w=1.66u
m10807 5522 5643 5500 VDDHV pch_18 l=0.27u w=1.66u
m10808 5523 5643 5501 VDDHV pch_18 l=0.27u w=1.66u
m10809 5524 5643 5502 VDDHV pch_18 l=0.27u w=1.66u
m10810 5551 5643 5535 VDDHV pch_18 l=0.27u w=1.66u
m10811 5552 5643 5536 VDDHV pch_18 l=0.27u w=1.66u
m10812 5553 5643 5537 VDDHV pch_18 l=0.27u w=1.66u
m10813 5554 5643 5538 VDDHV pch_18 l=0.27u w=1.66u
m10814 5555 5643 5539 VDDHV pch_18 l=0.27u w=1.66u
m10815 5556 5643 5540 VDDHV pch_18 l=0.27u w=1.66u
m10816 5557 5643 5541 VDDHV pch_18 l=0.27u w=1.66u
m10817 5558 5643 5542 VDDHV pch_18 l=0.27u w=1.66u
m10818 5559 5643 5543 VDDHV pch_18 l=0.27u w=1.66u
m10819 5560 5643 5544 VDDHV pch_18 l=0.27u w=1.66u
m10820 5561 5643 5545 VDDHV pch_18 l=0.27u w=1.66u
m10821 5562 5643 5546 VDDHV pch_18 l=0.27u w=1.66u
m10822 5582 5643 5567 VDDHV pch_18 l=0.27u w=1.66u
m10823 5583 5643 5568 VDDHV pch_18 l=0.27u w=1.66u
m10824 5584 5643 5569 VDDHV pch_18 l=0.27u w=1.66u
m10825 5585 5643 5570 VDDHV pch_18 l=0.27u w=1.66u
m10826 5586 5643 5571 VDDHV pch_18 l=0.27u w=1.66u
m10827 5587 5643 5572 VDDHV pch_18 l=0.27u w=1.66u
m10828 5588 5643 5573 VDDHV pch_18 l=0.27u w=1.66u
m10829 5589 5643 5574 VDDHV pch_18 l=0.27u w=1.66u
m10830 5590 5643 5575 VDDHV pch_18 l=0.27u w=1.66u
m10831 5591 5643 5576 VDDHV pch_18 l=0.27u w=1.66u
m10832 5592 5643 5577 VDDHV pch_18 l=0.27u w=1.66u
m10833 5593 5643 5578 VDDHV pch_18 l=0.27u w=1.66u
m10834 5067 5360 5506 VDDHV pch_18 l=0.28u w=0.44u
m10835 5615 5643 5598 VDDHV pch_18 l=0.27u w=1.66u
m10836 5616 5643 5599 VDDHV pch_18 l=0.27u w=1.66u
m10837 5617 5643 5600 VDDHV pch_18 l=0.27u w=1.66u
m10838 5618 5643 5601 VDDHV pch_18 l=0.27u w=1.66u
m10839 5619 5643 5602 VDDHV pch_18 l=0.27u w=1.66u
m10840 5620 5643 5603 VDDHV pch_18 l=0.27u w=1.66u
m10841 5621 5643 5604 VDDHV pch_18 l=0.27u w=1.66u
m10842 5622 5643 5605 VDDHV pch_18 l=0.27u w=1.66u
m10843 5623 5643 5606 VDDHV pch_18 l=0.27u w=1.66u
m10844 5624 5643 5607 VDDHV pch_18 l=0.27u w=1.66u
m10845 5625 5643 5608 VDDHV pch_18 l=0.27u w=1.66u
m10846 5626 5643 5609 VDDHV pch_18 l=0.27u w=1.66u
m10847 5645 5643 5631 VDDHV pch_18 l=0.27u w=1.66u
m10848 5646 5643 5632 VDDHV pch_18 l=0.27u w=1.66u
m10849 5647 5643 5633 VDDHV pch_18 l=0.27u w=1.66u
m10850 5648 5643 5634 VDDHV pch_18 l=0.27u w=1.66u
m10851 5649 5643 5635 VDDHV pch_18 l=0.27u w=1.66u
m10852 5650 5643 5636 VDDHV pch_18 l=0.27u w=1.66u
m10853 5651 5643 5637 VDDHV pch_18 l=0.27u w=1.66u
m10854 5652 5643 5638 VDDHV pch_18 l=0.27u w=1.66u
m10855 5653 5643 5639 VDDHV pch_18 l=0.27u w=1.66u
m10856 5654 5643 5640 VDDHV pch_18 l=0.27u w=1.66u
m10857 5655 5643 5641 VDDHV pch_18 l=0.27u w=1.66u
m10858 5656 5643 5642 VDDHV pch_18 l=0.27u w=1.66u
m10859 5677 5643 5663 VDDHV pch_18 l=0.27u w=1.66u
m10860 5678 5643 5664 VDDHV pch_18 l=0.27u w=1.66u
m10861 5679 5643 5665 VDDHV pch_18 l=0.27u w=1.66u
m10862 5680 5643 5666 VDDHV pch_18 l=0.27u w=1.66u
m10863 5681 5643 5667 VDDHV pch_18 l=0.27u w=1.66u
m10864 5682 5643 5668 VDDHV pch_18 l=0.27u w=1.66u
m10865 5683 5643 5669 VDDHV pch_18 l=0.27u w=1.66u
m10866 5684 5643 5670 VDDHV pch_18 l=0.27u w=1.66u
m10867 5685 5643 5671 VDDHV pch_18 l=0.27u w=1.66u
m10868 5686 5643 5672 VDDHV pch_18 l=0.27u w=1.66u
m10869 5687 5643 5673 VDDHV pch_18 l=0.27u w=1.66u
m10870 5688 5643 5674 VDDHV pch_18 l=0.27u w=1.66u
m10871 5709 5643 5694 VDDHV pch_18 l=0.27u w=1.66u
m10872 5710 5643 5695 VDDHV pch_18 l=0.27u w=1.66u
m10873 5711 5643 5696 VDDHV pch_18 l=0.27u w=1.66u
m10874 5712 5643 5697 VDDHV pch_18 l=0.27u w=1.66u
m10875 5713 5643 5698 VDDHV pch_18 l=0.27u w=1.66u
m10876 5714 5643 5699 VDDHV pch_18 l=0.27u w=1.66u
m10877 5715 5643 5700 VDDHV pch_18 l=0.27u w=1.66u
m10878 5716 5643 5701 VDDHV pch_18 l=0.27u w=1.66u
m10879 5717 5643 5702 VDDHV pch_18 l=0.27u w=1.66u
m10880 5718 5643 5703 VDDHV pch_18 l=0.27u w=1.66u
m10881 5719 5643 5704 VDDHV pch_18 l=0.27u w=1.66u
m10882 5720 5643 5705 VDDHV pch_18 l=0.27u w=1.66u
m10883 5726 5314 5067 VDDHV pch_18 l=0.28u w=0.44u
m10884 5734 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10885 5735 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10886 5736 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10887 5737 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10888 5738 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10889 5739 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10890 5740 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10891 5741 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10892 5742 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10893 5743 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10894 5744 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10895 5745 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10896 5753 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10897 5754 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10898 5755 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10899 5756 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10900 5757 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10901 5758 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10902 5759 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10903 5760 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10904 5761 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10905 5762 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10906 5763 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10907 5764 5643 5014 VDDHV pch_18 l=0.27u w=1.66u
m10908 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10909 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10910 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10911 5774 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10912 5775 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10913 5776 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10914 5777 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10915 5778 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10916 5779 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10917 5780 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10918 5781 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10919 5782 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10920 5786 5360 5726 VDDHV pch_18 l=0.28u w=0.44u
m10921 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10922 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10923 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10924 5774 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10925 5775 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10926 5776 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10927 5777 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10928 5778 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10929 5779 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10930 5780 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10931 5781 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10932 5782 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10933 VDDHV 5643 VDDHV VDDHV pch_18 l=0.27u w=1.66u
m10934 5803 5643 4994 VDDHV pch_18 l=0.27u w=1.66u
m10935 5804 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10936 5774 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10937 5775 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10938 5776 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10939 5777 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10940 5778 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10941 5779 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10942 5780 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10943 5781 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10944 5782 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10945 5815 5643 5809 VDDHV pch_18 l=0.27u w=1.66u
m10946 5816 5643 5786 VDDHV pch_18 l=0.27u w=1.66u
m10947 5804 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10948 5774 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10949 5775 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10950 5776 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10951 5777 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10952 5778 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10953 5779 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10954 5780 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10955 5781 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10956 5782 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10957 5830 5643 5784 VDDHV pch_18 l=0.27u w=1.66u
m10958 5816 5643 5786 VDDHV pch_18 l=0.27u w=1.66u
m10959 5804 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10960 5774 5643 5067 VDDHV pch_18 l=0.27u w=1.66u
m10961 5775 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10962 5776 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10963 5777 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10964 5778 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10965 5779 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10966 5780 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10967 5781 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10968 5782 5643 4 VDDHV pch_18 l=0.27u w=1.66u
m10969 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10970 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10971 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10972 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10973 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10974 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10975 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10976 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10977 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10978 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10979 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10980 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10981 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10982 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10983 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10984 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10985 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10986 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10987 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10988 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10989 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10990 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10991 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10992 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10993 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10994 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10995 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10996 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10997 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10998 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m10999 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11000 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11001 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11002 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11003 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11004 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11005 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11006 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11007 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11008 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11009 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11010 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11011 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11012 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11013 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11014 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11015 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11016 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11017 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11018 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11019 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11020 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11021 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11022 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11023 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11024 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11025 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11026 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11027 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11028 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11029 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11030 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11031 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11032 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11033 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11034 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11035 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11036 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11037 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11038 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11039 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11040 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11041 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11042 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11043 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11044 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11045 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11046 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11047 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11048 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11049 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11050 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11051 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11052 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11053 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11054 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11055 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11056 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11057 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11058 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11059 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11060 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11061 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11062 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11063 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11064 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11065 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11066 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11067 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11068 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11069 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11070 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11071 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11072 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11073 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11074 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11075 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11076 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11077 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11078 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11079 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11080 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11081 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11082 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11083 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11084 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11085 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11086 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11087 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11088 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11089 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11090 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11091 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11092 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11093 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11094 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11095 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11096 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11097 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11098 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11099 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11100 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11101 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11102 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11103 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11104 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11105 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11106 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11107 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11108 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11109 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11110 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11111 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11112 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11113 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11114 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11115 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11116 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11117 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11118 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11119 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11120 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11121 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11122 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11123 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11124 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11125 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11126 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11127 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11128 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11129 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11130 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11131 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11132 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11133 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11134 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11135 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11136 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11137 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11138 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11139 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11140 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11141 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11142 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11143 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11144 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11145 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11146 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11147 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11148 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11149 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11150 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11151 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11152 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11153 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11154 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11155 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11156 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11157 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11158 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11159 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11160 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11161 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11162 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11163 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11164 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11165 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11166 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11167 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11168 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11169 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11170 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11171 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11172 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11173 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11174 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11175 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11176 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11177 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11178 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11179 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11180 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11181 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11182 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11183 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11184 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11185 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11186 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11187 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11188 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11189 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11190 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11191 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11192 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11193 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11194 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11195 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11196 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11197 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11198 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11199 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11200 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11201 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11202 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11203 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11204 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11205 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11206 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11207 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11208 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11209 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11210 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11211 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11212 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11213 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11214 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11215 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11216 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11217 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11218 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11219 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11220 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11221 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11222 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11223 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11224 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11225 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11226 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11227 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11228 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11229 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11230 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11231 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11232 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11233 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11234 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11235 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11236 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11237 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11238 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11239 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11240 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11241 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11242 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11243 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11244 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11245 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11246 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11247 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11248 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11249 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11250 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11251 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11252 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11253 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11254 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11255 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11256 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11257 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11258 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11259 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11260 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11261 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11262 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11263 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11264 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11265 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11266 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11267 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11268 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11269 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11270 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11271 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11272 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11273 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11274 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11275 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11276 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11277 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11278 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11279 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11280 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11281 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11282 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11283 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11284 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11285 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11286 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11287 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11288 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11289 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11290 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11291 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11292 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11293 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11294 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11295 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11296 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11297 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11298 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11299 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11300 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11301 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11302 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11303 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11304 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11305 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11306 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11307 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11308 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11309 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11310 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11311 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11312 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11313 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11314 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11315 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11316 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11317 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11318 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11319 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11320 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11321 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11322 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11323 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11324 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11325 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11326 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11327 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11328 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11329 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11330 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11331 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11332 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11333 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11334 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11335 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11336 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11337 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11338 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11339 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11340 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11341 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11342 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11343 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11344 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11345 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11346 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11347 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11348 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11349 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11350 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11351 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11352 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11353 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11354 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11355 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11356 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11357 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11358 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11359 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11360 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11361 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11362 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11363 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11364 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11365 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11366 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11367 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11368 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11369 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11370 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11371 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11372 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11373 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11374 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11375 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11376 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11377 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11378 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11379 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11380 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11381 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11382 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11383 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11384 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11385 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11386 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11387 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11388 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11389 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11390 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11391 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11392 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11393 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11394 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11395 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11396 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11397 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11398 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11399 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11400 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11401 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11402 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11403 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11404 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11405 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11406 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11407 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11408 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11409 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11410 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11411 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11412 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11413 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11414 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11415 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11416 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11417 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11418 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11419 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11420 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11421 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11422 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11423 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11424 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11425 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11426 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11427 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11428 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11429 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11430 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11431 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11432 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11433 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11434 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11435 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11436 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11437 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11438 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11439 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11440 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11441 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11442 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11443 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11444 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11445 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11446 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11447 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11448 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11449 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11450 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11451 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11452 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11453 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11454 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11455 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11456 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11457 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11458 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11459 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11460 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11461 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11462 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11463 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11464 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11465 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11466 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11467 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11468 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11469 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11470 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11471 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11472 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11473 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11474 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11475 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11476 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11477 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11478 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11479 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11480 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11481 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11482 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11483 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11484 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11485 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11486 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11487 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11488 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11489 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11490 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11491 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11492 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11493 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11494 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11495 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11496 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11497 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11498 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11499 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11500 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11501 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11502 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11503 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11504 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11505 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11506 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11507 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11508 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11509 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11510 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11511 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11512 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11513 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11514 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11515 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11516 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11517 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11518 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11519 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11520 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11521 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11522 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11523 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11524 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11525 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11526 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11527 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11528 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11529 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11530 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11531 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11532 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11533 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11534 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11535 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11536 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11537 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11538 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11539 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11540 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11541 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11542 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11543 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11544 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11545 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11546 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11547 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11548 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11549 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11550 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11551 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11552 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11553 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11554 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11555 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11556 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11557 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11558 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11559 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11560 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11561 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11562 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11563 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11564 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11565 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11566 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11567 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11568 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11569 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11570 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11571 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11572 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11573 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11574 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11575 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11576 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11577 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11578 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11579 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11580 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11581 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11582 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11583 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11584 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11585 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11586 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11587 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11588 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11589 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11590 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11591 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11592 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11593 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11594 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11595 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11596 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11597 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11598 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11599 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11600 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11601 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11602 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11603 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11604 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11605 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11606 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11607 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11608 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11609 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11610 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11611 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11612 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11613 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11614 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11615 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11616 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11617 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11618 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11619 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11620 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11621 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11622 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11623 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11624 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11625 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11626 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11627 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11628 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11629 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11630 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11631 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11632 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11633 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11634 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11635 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11636 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11637 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11638 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11639 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11640 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11641 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11642 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11643 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11644 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11645 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11646 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11647 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11648 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11649 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11650 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11651 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11652 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11653 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11654 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11655 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11656 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11657 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11658 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11659 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11660 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11661 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11662 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11663 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11664 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11665 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11666 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11667 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11668 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11669 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11670 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11671 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11672 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11673 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11674 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11675 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11676 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11677 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11678 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11679 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11680 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11681 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11682 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11683 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11684 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11685 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11686 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11687 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11688 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11689 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11690 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11691 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11692 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11693 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11694 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11695 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11696 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11697 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11698 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11699 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11700 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11701 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11702 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11703 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11704 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11705 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11706 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11707 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11708 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11709 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11710 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11711 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11712 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11713 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11714 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11715 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11716 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11717 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11718 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11719 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11720 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11721 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11722 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11723 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11724 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11725 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11726 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11727 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11728 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11729 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11730 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11731 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11732 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11733 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11734 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11735 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11736 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11737 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11738 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11739 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11740 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11741 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11742 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11743 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11744 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11745 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11746 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11747 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11748 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11749 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11750 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11751 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11752 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11753 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11754 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11755 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11756 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11757 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11758 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11759 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11760 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11761 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11762 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11763 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11764 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11765 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11766 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11767 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11768 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11769 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11770 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11771 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11772 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11773 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11774 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11775 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11776 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11777 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11778 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11779 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11780 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11781 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11782 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11783 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11784 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11785 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11786 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11787 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11788 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11789 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11790 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11791 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11792 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11793 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11794 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11795 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11796 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11797 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11798 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11799 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11800 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11801 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11802 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11803 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11804 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11805 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11806 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11807 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11808 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11809 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11810 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11811 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11812 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11813 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11814 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11815 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11816 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11817 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11818 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11819 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11820 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11821 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11822 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11823 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11824 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11825 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11826 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11827 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11828 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11829 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11830 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11831 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11832 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11833 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11834 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11835 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11836 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11837 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11838 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11839 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11840 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11841 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11842 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11843 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11844 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11845 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11846 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11847 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11848 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11849 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11850 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11851 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11852 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11853 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11854 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11855 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11856 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11857 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11858 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11859 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11860 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11861 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11862 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11863 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11864 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11865 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11866 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11867 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11868 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11869 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11870 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11871 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11872 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11873 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11874 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11875 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11876 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11877 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11878 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11879 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11880 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11881 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11882 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11883 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11884 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11885 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11886 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11887 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11888 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11889 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11890 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11891 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11892 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11893 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11894 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11895 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11896 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11897 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11898 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11899 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11900 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11901 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11902 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11903 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11904 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11905 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11906 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11907 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11908 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11909 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11910 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11911 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11912 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11913 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11914 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11915 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11916 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11917 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11918 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11919 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11920 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11921 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11922 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11923 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11924 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11925 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11926 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11927 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11928 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11929 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11930 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11931 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11932 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11933 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11934 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11935 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11936 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11937 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11938 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11939 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11940 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11941 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11942 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11943 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11944 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11945 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11946 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11947 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11948 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11949 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11950 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11951 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11952 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11953 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11954 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11955 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11956 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11957 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11958 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11959 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11960 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11961 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11962 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11963 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11964 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11965 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11966 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11967 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11968 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11969 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11970 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11971 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11972 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11973 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11974 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11975 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11976 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11977 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11978 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11979 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11980 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11981 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11982 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11983 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11984 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11985 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11986 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11987 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11988 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11989 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11990 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11991 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11992 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11993 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11994 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11995 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11996 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11997 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11998 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m11999 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12000 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12001 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12002 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12003 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12004 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12005 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12006 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12007 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12008 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12009 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12010 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12011 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12012 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12013 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12014 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12015 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12016 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12017 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12018 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12019 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12020 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12021 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12022 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12023 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12024 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12025 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12026 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12027 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12028 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12029 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12030 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12031 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12032 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12033 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12034 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12035 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12036 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12037 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12038 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12039 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12040 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12041 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12042 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12043 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12044 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12045 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12046 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12047 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12048 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12049 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12050 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12051 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12052 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12053 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12054 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12055 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12056 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12057 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12058 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12059 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12060 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12061 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12062 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12063 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12064 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12065 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12066 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12067 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12068 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12069 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12070 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12071 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12072 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12073 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12074 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12075 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12076 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12077 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12078 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12079 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12080 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12081 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12082 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12083 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12084 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12085 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12086 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12087 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12088 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12089 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12090 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12091 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12092 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12093 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12094 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12095 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12096 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12097 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12098 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12099 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12100 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12101 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12102 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12103 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12104 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12105 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12106 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12107 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12108 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12109 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12110 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12111 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12112 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12113 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12114 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12115 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12116 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12117 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12118 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12119 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12120 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12121 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12122 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12123 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12124 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12125 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12126 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12127 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12128 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12129 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12130 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12131 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12132 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12133 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12134 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12135 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12136 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12137 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12138 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12139 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12140 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12141 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12142 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12143 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12144 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12145 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12146 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12147 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12148 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12149 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12150 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12151 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12152 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12153 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12154 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12155 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12156 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12157 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12158 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12159 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12160 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12161 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12162 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12163 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12164 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12165 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12166 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12167 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12168 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12169 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12170 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12171 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12172 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12173 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12174 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12175 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12176 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12177 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12178 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12179 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12180 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12181 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12182 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12183 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12184 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12185 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12186 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12187 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12188 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12189 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12190 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12191 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12192 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12193 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12194 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12195 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12196 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12197 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12198 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12199 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12200 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12201 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12202 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12203 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12204 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12205 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12206 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12207 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12208 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12209 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12210 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12211 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12212 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12213 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12214 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12215 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12216 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12217 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12218 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12219 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12220 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12221 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12222 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12223 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12224 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12225 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12226 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12227 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12228 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12229 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12230 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12231 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12232 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12233 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12234 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12235 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12236 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12237 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12238 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12239 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12240 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12241 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12242 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12243 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12244 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12245 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12246 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12247 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12248 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12249 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12250 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12251 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12252 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12253 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12254 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12255 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12256 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12257 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12258 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12259 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12260 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12261 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12262 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12263 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12264 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12265 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12266 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12267 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12268 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12269 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12270 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12271 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12272 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12273 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12274 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12275 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12276 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12277 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12278 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12279 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12280 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12281 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12282 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12283 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12284 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12285 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12286 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12287 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12288 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12289 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12290 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12291 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12292 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12293 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12294 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12295 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12296 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12297 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12298 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12299 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12300 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12301 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12302 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12303 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12304 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12305 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12306 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12307 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12308 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12309 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12310 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12311 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12312 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12313 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12314 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12315 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12316 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12317 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12318 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12319 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12320 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12321 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12322 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12323 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12324 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12325 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12326 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12327 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12328 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12329 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12330 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12331 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12332 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12333 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12334 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12335 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12336 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12337 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12338 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12339 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12340 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12341 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12342 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12343 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12344 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12345 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12346 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12347 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12348 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12349 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12350 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12351 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12352 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12353 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12354 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12355 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12356 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12357 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12358 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12359 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12360 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12361 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12362 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12363 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12364 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12365 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12366 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12367 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12368 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12369 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12370 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12371 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12372 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12373 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12374 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12375 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12376 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12377 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12378 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12379 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12380 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12381 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12382 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12383 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12384 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12385 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12386 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12387 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12388 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12389 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12390 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12391 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12392 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12393 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12394 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12395 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12396 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12397 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12398 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12399 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12400 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12401 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12402 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12403 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12404 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12405 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12406 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12407 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12408 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12409 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12410 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12411 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12412 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12413 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12414 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12415 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12416 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12417 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12418 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12419 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12420 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12421 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12422 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12423 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12424 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12425 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12426 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12427 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12428 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12429 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12430 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12431 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12432 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12433 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12434 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12435 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12436 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12437 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12438 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12439 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12440 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12441 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12442 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12443 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12444 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12445 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12446 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12447 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12448 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12449 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12450 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12451 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12452 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12453 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12454 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12455 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12456 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12457 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12458 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12459 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12460 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12461 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12462 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12463 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12464 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12465 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12466 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12467 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12468 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12469 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12470 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12471 VDDHV 2 4717 VDDHV pch_18 l=0.65u w=0.975u
m12472 4718 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12473 VDDHV 2 4719 VDDHV pch_18 l=0.65u w=0.975u
m12474 4720 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12475 VDDHV 2 4721 VDDHV pch_18 l=0.65u w=0.975u
m12476 4722 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12477 VDDHV 2 4723 VDDHV pch_18 l=0.65u w=0.975u
m12478 4724 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12479 VDDHV 2 4725 VDDHV pch_18 l=0.65u w=0.975u
m12480 4726 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12481 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12482 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12483 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12484 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12485 VDDHV 2 4727 VDDHV pch_18 l=0.65u w=0.975u
m12486 4728 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12487 VDDHV 2 4729 VDDHV pch_18 l=0.65u w=0.975u
m12488 4730 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12489 VDDHV 2 4731 VDDHV pch_18 l=0.65u w=0.975u
m12490 4732 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12491 VDDHV 2 4733 VDDHV pch_18 l=0.65u w=0.975u
m12492 4734 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12493 VDDHV 2 4735 VDDHV pch_18 l=0.65u w=0.975u
m12494 4736 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12495 VDDHV 2 4737 VDDHV pch_18 l=0.65u w=0.975u
m12496 4737 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12497 VDDHV 2 4738 VDDHV pch_18 l=0.65u w=0.975u
m12498 4738 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12499 VDDHV 2 4739 VDDHV pch_18 l=0.65u w=0.975u
m12500 4740 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12501 VDDHV 2 4741 VDDHV pch_18 l=0.65u w=0.975u
m12502 4742 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12503 VDDHV 2 4743 VDDHV pch_18 l=0.65u w=0.975u
m12504 4744 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12505 VDDHV 2 4745 VDDHV pch_18 l=0.65u w=0.975u
m12506 4746 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12507 VDDHV 2 4747 VDDHV pch_18 l=0.65u w=0.975u
m12508 4748 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12509 VDDHV 2 4749 VDDHV pch_18 l=0.65u w=0.975u
m12510 4749 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12511 VDDHV 2 4750 VDDHV pch_18 l=0.65u w=0.975u
m12512 4750 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12513 VDDHV 2 4751 VDDHV pch_18 l=0.65u w=0.975u
m12514 4752 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12515 VDDHV 2 4753 VDDHV pch_18 l=0.65u w=0.975u
m12516 4754 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12517 VDDHV 2 4755 VDDHV pch_18 l=0.65u w=0.975u
m12518 4756 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12519 VDDHV 2 4757 VDDHV pch_18 l=0.65u w=0.975u
m12520 4758 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12521 VDDHV 2 4759 VDDHV pch_18 l=0.65u w=0.975u
m12522 4760 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12523 VDDHV 2 4761 VDDHV pch_18 l=0.65u w=0.975u
m12524 4761 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12525 VDDHV 2 4762 VDDHV pch_18 l=0.65u w=0.975u
m12526 4762 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12527 VDDHV 2 4763 VDDHV pch_18 l=0.65u w=0.975u
m12528 4764 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12529 VDDHV 2 4765 VDDHV pch_18 l=0.65u w=0.975u
m12530 4766 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12531 VDDHV 2 4767 VDDHV pch_18 l=0.65u w=0.975u
m12532 4768 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12533 VDDHV 2 4769 VDDHV pch_18 l=0.65u w=0.975u
m12534 4770 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12535 VDDHV 2 4771 VDDHV pch_18 l=0.65u w=0.975u
m12536 4772 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12537 VDDHV 2 4773 VDDHV pch_18 l=0.65u w=0.975u
m12538 4773 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12539 VDDHV 2 4774 VDDHV pch_18 l=0.65u w=0.975u
m12540 4774 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12541 VDDHV 2 4775 VDDHV pch_18 l=0.65u w=0.975u
m12542 4776 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12543 VDDHV 2 4777 VDDHV pch_18 l=0.65u w=0.975u
m12544 4778 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12545 VDDHV 2 4779 VDDHV pch_18 l=0.65u w=0.975u
m12546 4780 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12547 VDDHV 2 4781 VDDHV pch_18 l=0.65u w=0.975u
m12548 4782 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12549 VDDHV 2 4783 VDDHV pch_18 l=0.65u w=0.975u
m12550 4784 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12551 VDDHV 2 4785 VDDHV pch_18 l=0.65u w=0.975u
m12552 4785 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12553 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12554 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12555 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12556 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12557 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12558 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12559 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12560 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12561 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12562 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12563 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12564 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12565 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12566 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12567 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12568 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12569 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12570 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12571 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12572 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12573 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12574 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12575 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12576 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12577 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12578 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12579 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12580 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12581 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12582 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12583 4859 VSS VDDHV VDDHV pch_18 l=10u w=0.44u
m12584 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12585 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12586 VDDHV 2 4797 VDDHV pch_18 l=0.65u w=0.975u
m12587 4798 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12588 VDDHV 2 4799 VDDHV pch_18 l=0.65u w=0.975u
m12589 4800 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12590 VDDHV 2 4801 VDDHV pch_18 l=0.65u w=0.975u
m12591 4802 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12592 VDDHV 2 4803 VDDHV pch_18 l=0.65u w=0.975u
m12593 4804 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12594 VDDHV 2 4805 VDDHV pch_18 l=0.65u w=0.975u
m12595 4806 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12596 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12597 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12598 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12599 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12600 VDDHV 2 4807 VDDHV pch_18 l=0.65u w=0.975u
m12601 4808 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12602 VDDHV 2 4809 VDDHV pch_18 l=0.65u w=0.975u
m12603 4810 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12604 VDDHV 2 4811 VDDHV pch_18 l=0.65u w=0.975u
m12605 4812 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12606 VDDHV 2 4813 VDDHV pch_18 l=0.65u w=0.975u
m12607 4814 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12608 VDDHV 2 4815 VDDHV pch_18 l=0.65u w=0.975u
m12609 4816 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12610 VDDHV 2 4737 VDDHV pch_18 l=0.65u w=0.975u
m12611 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12612 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12613 4738 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12614 VDDHV 2 4817 VDDHV pch_18 l=0.65u w=0.975u
m12615 4818 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12616 VDDHV 2 4819 VDDHV pch_18 l=0.65u w=0.975u
m12617 4820 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12618 VDDHV 2 4821 VDDHV pch_18 l=0.65u w=0.975u
m12619 4822 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12620 VDDHV 2 4823 VDDHV pch_18 l=0.65u w=0.975u
m12621 4824 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12622 VDDHV 2 4825 VDDHV pch_18 l=0.65u w=0.975u
m12623 4826 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12624 VDDHV 2 4749 VDDHV pch_18 l=0.65u w=0.975u
m12625 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12626 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12627 4750 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12628 VDDHV 2 4827 VDDHV pch_18 l=0.65u w=0.975u
m12629 4828 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12630 VDDHV 2 4829 VDDHV pch_18 l=0.65u w=0.975u
m12631 4830 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12632 VDDHV 2 4831 VDDHV pch_18 l=0.65u w=0.975u
m12633 4832 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12634 VDDHV 2 4833 VDDHV pch_18 l=0.65u w=0.975u
m12635 4834 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12636 VDDHV 2 4835 VDDHV pch_18 l=0.65u w=0.975u
m12637 4836 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12638 VDDHV 2 4761 VDDHV pch_18 l=0.65u w=0.975u
m12639 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12640 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12641 4762 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12642 VDDHV 2 4837 VDDHV pch_18 l=0.65u w=0.975u
m12643 4838 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12644 VDDHV 2 4839 VDDHV pch_18 l=0.65u w=0.975u
m12645 4840 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12646 VDDHV 2 4841 VDDHV pch_18 l=0.65u w=0.975u
m12647 4842 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12648 VDDHV 2 4843 VDDHV pch_18 l=0.65u w=0.975u
m12649 4844 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12650 VDDHV 2 4845 VDDHV pch_18 l=0.65u w=0.975u
m12651 4846 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12652 VDDHV 2 4773 VDDHV pch_18 l=0.65u w=0.975u
m12653 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12654 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12655 4774 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12656 VDDHV 2 4847 VDDHV pch_18 l=0.65u w=0.975u
m12657 4848 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12658 VDDHV 2 4849 VDDHV pch_18 l=0.65u w=0.975u
m12659 4850 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12660 VDDHV 2 4851 VDDHV pch_18 l=0.65u w=0.975u
m12661 4852 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12662 VDDHV 2 4853 VDDHV pch_18 l=0.65u w=0.975u
m12663 4854 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12664 VDDHV 2 4855 VDDHV pch_18 l=0.65u w=0.975u
m12665 4856 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12666 VDDHV 2 4785 VDDHV pch_18 l=0.65u w=0.975u
m12667 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12668 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12669 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12670 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12671 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12672 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12673 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12674 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12675 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12676 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12677 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12678 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12679 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12680 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12681 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12682 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12683 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12684 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12685 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12686 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12687 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12688 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12689 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12690 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12691 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12692 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12693 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12694 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12695 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12696 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12697 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12698 4868 4795 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12699 4869 4949 4868 VDDHV pch_18 l=0.44u w=1.04u
m12700 VDDHV 4859 4865 VDDHV pch_18 l=0.44u w=1.04u
m12701 4864 4869 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12702 VDDHV 4795 4796 VDDHV pch_18 l=0.44u w=1.04u
m12703 4795 4948 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12704 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12705 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12706 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12707 4877 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12708 VDDHV 2 4878 VDDHV pch_18 l=0.65u w=0.975u
m12709 4879 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12710 VDDHV 2 4880 VDDHV pch_18 l=0.65u w=0.975u
m12711 4881 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12712 VDDHV 2 4882 VDDHV pch_18 l=0.65u w=0.975u
m12713 4883 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12714 VDDHV 2 4884 VDDHV pch_18 l=0.65u w=0.975u
m12715 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12716 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12717 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12718 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12719 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12720 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12721 4885 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12722 VDDHV 2 4886 VDDHV pch_18 l=0.65u w=0.975u
m12723 4887 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12724 VDDHV 2 4888 VDDHV pch_18 l=0.65u w=0.975u
m12725 4889 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12726 VDDHV 2 4890 VDDHV pch_18 l=0.65u w=0.975u
m12727 4891 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12728 VDDHV 2 4892 VDDHV pch_18 l=0.65u w=0.975u
m12729 4737 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12730 VDDHV 2 4737 VDDHV pch_18 l=0.65u w=0.975u
m12731 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12732 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12733 4738 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12734 VDDHV 2 4738 VDDHV pch_18 l=0.65u w=0.975u
m12735 4893 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12736 VDDHV 2 4894 VDDHV pch_18 l=0.65u w=0.975u
m12737 4895 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12738 VDDHV 2 4896 VDDHV pch_18 l=0.65u w=0.975u
m12739 4897 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12740 VDDHV 2 4898 VDDHV pch_18 l=0.65u w=0.975u
m12741 4899 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12742 VDDHV 2 4900 VDDHV pch_18 l=0.65u w=0.975u
m12743 4749 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12744 VDDHV 2 4749 VDDHV pch_18 l=0.65u w=0.975u
m12745 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12746 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12747 4750 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12748 VDDHV 2 4750 VDDHV pch_18 l=0.65u w=0.975u
m12749 4901 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12750 VDDHV 2 4902 VDDHV pch_18 l=0.65u w=0.975u
m12751 4903 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12752 VDDHV 2 4904 VDDHV pch_18 l=0.65u w=0.975u
m12753 4905 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12754 VDDHV 2 4906 VDDHV pch_18 l=0.65u w=0.975u
m12755 4907 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12756 VDDHV 2 4908 VDDHV pch_18 l=0.65u w=0.975u
m12757 4761 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12758 VDDHV 2 4761 VDDHV pch_18 l=0.65u w=0.975u
m12759 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12760 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12761 4762 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12762 VDDHV 2 4762 VDDHV pch_18 l=0.65u w=0.975u
m12763 4909 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12764 VDDHV 2 4910 VDDHV pch_18 l=0.65u w=0.975u
m12765 4911 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12766 VDDHV 2 4912 VDDHV pch_18 l=0.65u w=0.975u
m12767 4913 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12768 VDDHV 2 4914 VDDHV pch_18 l=0.65u w=0.975u
m12769 4915 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12770 VDDHV 2 4916 VDDHV pch_18 l=0.65u w=0.975u
m12771 4773 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12772 VDDHV 2 4773 VDDHV pch_18 l=0.65u w=0.975u
m12773 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12774 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12775 4774 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12776 VDDHV 2 4774 VDDHV pch_18 l=0.65u w=0.975u
m12777 4917 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12778 VDDHV 2 4918 VDDHV pch_18 l=0.65u w=0.975u
m12779 4919 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12780 VDDHV 2 4920 VDDHV pch_18 l=0.65u w=0.975u
m12781 4921 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12782 VDDHV 2 4922 VDDHV pch_18 l=0.65u w=0.975u
m12783 4923 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12784 VDDHV 2 4924 VDDHV pch_18 l=0.65u w=0.975u
m12785 4785 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12786 VDDHV 2 4785 VDDHV pch_18 l=0.65u w=0.975u
m12787 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m12788 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12789 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12790 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12791 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12792 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12793 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12794 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12795 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12796 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12797 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12798 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12799 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12800 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12801 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12802 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12803 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12804 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12805 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12806 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12807 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12808 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12809 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12810 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12811 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12812 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12813 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12814 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12815 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12816 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12817 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12818 42575 4938 VDDHV VDDHV pch_18 l=0.8u w=0.44u
m12819 42576 4938 42575 VDDHV pch_18 l=0.8u w=0.44u
m12820 42577 4938 42576 VDDHV pch_18 l=0.8u w=0.44u
m12821 42578 4938 42577 VDDHV pch_18 l=0.8u w=0.44u
m12822 4859 4946 42578 VDDHV pch_18 l=0.44u w=0.44u
m12823 VDDHV 4865 2 VDDHV pch_18 l=1.04u w=2.08u
m12824 4948 VSS 4867 VDDHV pch_18 l=4.5u w=0.44u
m12825 VDDHV VSS 4867 VDDHV pch_18 l=4.5u w=0.44u
m12826 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12827 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12828 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12829 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12830 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12831 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12832 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12833 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12834 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12835 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12836 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12837 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12838 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12839 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12840 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12841 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12842 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12843 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12844 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12845 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12846 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12847 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12848 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12849 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12850 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12851 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12852 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12853 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12854 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12855 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12856 43526 4938 VDDHV VDDHV pch_18 l=0.8u w=0.44u
m12857 43527 4938 43526 VDDHV pch_18 l=0.8u w=0.44u
m12858 43528 4938 43527 VDDHV pch_18 l=0.8u w=0.44u
m12859 43529 4938 43528 VDDHV pch_18 l=0.8u w=0.44u
m12860 4946 4859 43529 VDDHV pch_18 l=0.44u w=0.44u
m12861 43991 4957 VDDHV VDDHV pch_18 l=0.8u w=0.44u
m12862 43992 4957 43991 VDDHV pch_18 l=0.8u w=0.44u
m12863 43993 4957 43992 VDDHV pch_18 l=0.8u w=0.44u
m12864 43994 4957 43993 VDDHV pch_18 l=0.8u w=0.44u
m12865 4954 4948 43994 VDDHV pch_18 l=0.44u w=0.44u
m12866 4861 4796 2 VDDHV pch_18 l=0.44u w=2.08u
m12867 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12868 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12869 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12870 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12871 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12872 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12873 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12874 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12875 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12876 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12877 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12878 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12879 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12880 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12881 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12882 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12883 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12884 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12885 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12886 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12887 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12888 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12889 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12890 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12891 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12892 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12893 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12894 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12895 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12896 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12897 44470 4957 VDDHV VDDHV pch_18 l=0.8u w=0.44u
m12898 44471 4957 44470 VDDHV pch_18 l=0.8u w=0.44u
m12899 44472 4957 44471 VDDHV pch_18 l=0.8u w=0.44u
m12900 44473 4957 44472 VDDHV pch_18 l=0.8u w=0.44u
m12901 4948 4954 44473 VDDHV pch_18 l=0.44u w=0.44u
m12902 45178 4975 VDDHV VDDHV pch_18 l=0.8u w=0.44u
m12903 45179 4975 45178 VDDHV pch_18 l=0.8u w=0.44u
m12904 45180 4975 45179 VDDHV pch_18 l=0.8u w=0.44u
m12905 45181 4975 45180 VDDHV pch_18 l=0.8u w=0.44u
m12906 4971 4949 45181 VDDHV pch_18 l=0.44u w=0.44u
m12907 4862 4864 2 VDDHV pch_18 l=0.44u w=2.08u
m12908 4988 VSS 4949 VDDHV pch_18 l=4.5u w=0.44u
m12909 4988 VSS VDDHV VDDHV pch_18 l=4.5u w=0.44u
m12910 46404 4975 VDDHV VDDHV pch_18 l=0.8u w=0.44u
m12911 46405 4975 46404 VDDHV pch_18 l=0.8u w=0.44u
m12912 46406 4975 46405 VDDHV pch_18 l=0.8u w=0.44u
m12913 46407 4975 46406 VDDHV pch_18 l=0.8u w=0.44u
m12914 4949 4971 46407 VDDHV pch_18 l=0.44u w=0.44u
m12915 5001 5068 4992 VDDHV pch_18 l=0.44u w=1.04u
m12916 5001 5068 4992 VDDHV pch_18 l=0.44u w=1.04u
m12917 VDDHV 4992 4996 VDDHV pch_18 l=0.44u w=1.04u
m12918 47493 5068 4992 VDDHV pch_18 l=0.44u w=0.44u
m12919 VDDHV 5020 5001 VDDHV pch_18 l=0.44u w=1.04u
m12920 VDDHV 5020 5001 VDDHV pch_18 l=0.44u w=1.04u
m12921 5020 4996 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12922 5020 4996 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12923 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12924 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12925 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12926 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12927 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12928 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12929 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12930 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12931 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12932 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12933 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12934 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12935 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12936 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12937 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12938 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12939 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12940 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12941 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12942 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12943 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12944 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12945 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12946 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12947 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12948 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12949 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12950 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12951 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12952 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12953 5001 5020 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12954 5001 5020 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12955 VDDHV VSS 47493 VDDHV pch_18 l=0.8u w=0.44u
m12956 VDDHV 4996 5020 VDDHV pch_18 l=0.44u w=1.04u
m12957 VDDHV 4996 5020 VDDHV pch_18 l=0.44u w=1.04u
m12958 5048 5072 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12959 5048 5072 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12960 VDDHV 5048 5043 VDDHV pch_18 l=0.44u w=1.04u
m12961 VDDHV 5048 5043 VDDHV pch_18 l=0.44u w=1.04u
m12962 48193 VSS VDDHV VDDHV pch_18 l=0.8u w=0.44u
m12963 VDDHV 5072 5048 VDDHV pch_18 l=0.44u w=1.04u
m12964 VDDHV 5072 5048 VDDHV pch_18 l=0.44u w=1.04u
m12965 5043 5048 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12966 5043 5048 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12967 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12968 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12969 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12970 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12971 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12972 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12973 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12974 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12975 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12976 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12977 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12978 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12979 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12980 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12981 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12982 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12983 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12984 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12985 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12986 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12987 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12988 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12989 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12990 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12991 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12992 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12993 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12994 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12995 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12996 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m12997 5068 4992 48193 VDDHV pch_18 l=0.44u w=0.44u
m12998 5072 5068 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m12999 5068 4992 5043 VDDHV pch_18 l=0.44u w=1.04u
m13000 5068 4992 5043 VDDHV pch_18 l=0.44u w=1.04u
m13001 5068 VSS 4991 VDDHV pch_18 l=5u w=0.44u
m13002 VDDHV VSS 4991 VDDHV pch_18 l=5u w=0.44u
m13003 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13004 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13005 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13006 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13007 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13008 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13009 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13010 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13011 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13012 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13013 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13014 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13015 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13016 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13017 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13018 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13019 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13020 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13021 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13022 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13023 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13024 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13025 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13026 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13027 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13028 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13029 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13030 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13031 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13032 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13033 5114 5178 5093 VDDHV pch_18 l=0.44u w=1.04u
m13034 5114 5178 5093 VDDHV pch_18 l=0.44u w=1.04u
m13035 VDDHV 5093 5097 VDDHV pch_18 l=0.44u w=1.04u
m13036 49415 5178 5093 VDDHV pch_18 l=0.44u w=0.44u
m13037 VDDHV 5131 5114 VDDHV pch_18 l=0.44u w=1.04u
m13038 VDDHV 5131 5114 VDDHV pch_18 l=0.44u w=1.04u
m13039 5131 5097 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13040 5131 5097 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13041 5114 5131 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13042 5114 5131 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13043 VDDHV VSS 49415 VDDHV pch_18 l=0.8u w=0.44u
m13044 VDDHV 5097 5131 VDDHV pch_18 l=0.44u w=1.04u
m13045 VDDHV 5097 5131 VDDHV pch_18 l=0.44u w=1.04u
m13046 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13047 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13048 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13049 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13050 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13051 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13052 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13053 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13054 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13055 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13056 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13057 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13058 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13059 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13060 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13061 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13062 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13063 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13064 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13065 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13066 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13067 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13068 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13069 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13070 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13071 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13072 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13073 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13074 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13075 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13076 5158 5183 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13077 5158 5183 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13078 VDDHV 5158 5141 VDDHV pch_18 l=0.44u w=1.04u
m13079 VDDHV 5158 5141 VDDHV pch_18 l=0.44u w=1.04u
m13080 50054 VSS VDDHV VDDHV pch_18 l=0.8u w=0.44u
m13081 VDDHV 5183 5158 VDDHV pch_18 l=0.44u w=1.04u
m13082 VDDHV 5183 5158 VDDHV pch_18 l=0.44u w=1.04u
m13083 5141 5158 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13084 5141 5158 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13085 5178 5093 50054 VDDHV pch_18 l=0.44u w=0.44u
m13086 5183 5178 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13087 5178 5093 5141 VDDHV pch_18 l=0.44u w=1.04u
m13088 5178 5093 5141 VDDHV pch_18 l=0.44u w=1.04u
m13089 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13090 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13091 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13092 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13093 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13094 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13095 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13096 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13097 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13098 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13099 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13100 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13101 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13102 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13103 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13104 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13105 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13106 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13107 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13108 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13109 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13110 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13111 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13112 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13113 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13114 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13115 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13116 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13117 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13118 VDDHV 4862 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13119 5178 VSS 5092 VDDHV pch_18 l=5u w=0.44u
m13120 VDDHV VSS 5092 VDDHV pch_18 l=5u w=0.44u
m13121 VDDHV 5048 5205 VDDHV pch_18 l=0.44u w=1.04u
m13122 5231 5020 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13123 5234 5205 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13124 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13125 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13126 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13127 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13128 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13129 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13130 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13131 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13132 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13133 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13134 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13135 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13136 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13137 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13138 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13139 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13140 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13141 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13142 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13143 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13144 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13145 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13146 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13147 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13148 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13149 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13150 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13151 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13152 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13153 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13154 VDDHV 5273 5249 VDDHV pch_18 l=0.44u w=1.04u
m13155 VDDHV 5131 5250 VDDHV pch_18 l=0.44u w=1.04u
m13156 5273 5158 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13157 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13158 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13159 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13160 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13161 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13162 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13163 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13164 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13165 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13166 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13167 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13168 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13169 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13170 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13171 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13172 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13173 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13174 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13175 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13176 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13177 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13178 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13179 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13180 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13181 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13182 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13183 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13184 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13185 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13186 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13187 VDDHV VDDHV VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13188 VDDHV VDDHV VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13189 VDDHV VDDHV VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13190 VDDHV VDDHV VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13191 5316 5315 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13192 5313 5312 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13193 5315 5158 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13194 5312 5131 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13195 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13196 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13197 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13198 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13199 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13200 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13201 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13202 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13203 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13204 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13205 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13206 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13207 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13208 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13209 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13210 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13211 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13212 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13213 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13214 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13215 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13216 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13217 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13218 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13219 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13220 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13221 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13222 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13223 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13224 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13225 VDDHV 5315 5316 VDDHV pch_18 l=0.44u w=1.04u
m13226 VDDHV 5312 5313 VDDHV pch_18 l=0.44u w=1.04u
m13227 VDDHV 5158 5315 VDDHV pch_18 l=0.44u w=1.04u
m13228 VDDHV 5131 5312 VDDHV pch_18 l=0.44u w=1.04u
m13229 5356 5358 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13230 5357 5359 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13231 5358 5048 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13232 5359 5020 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13233 VDDHV 5358 5356 VDDHV pch_18 l=0.44u w=1.04u
m13234 VDDHV 5359 5357 VDDHV pch_18 l=0.44u w=1.04u
m13235 VDDHV 5048 5358 VDDHV pch_18 l=0.44u w=1.04u
m13236 VDDHV 5020 5359 VDDHV pch_18 l=0.44u w=1.04u
m13237 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13238 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13239 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13240 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13241 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13242 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13243 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13244 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13245 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13246 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13247 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13248 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13249 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13250 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13251 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13252 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13253 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13254 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13255 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13256 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13257 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13258 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13259 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13260 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13261 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13262 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13263 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13264 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13265 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13266 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13267 5314 5357 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13268 5314 5357 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13269 5360 5356 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13270 5360 5356 VDDHV VDDHV pch_18 l=0.44u w=1.04u
m13271 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13272 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13273 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13274 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13275 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13276 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13277 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13278 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13279 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13280 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13281 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13282 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13283 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13284 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13285 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13286 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13287 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13288 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13289 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13290 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13291 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13292 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13293 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13294 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13295 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13296 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13297 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13298 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13299 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13300 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13301 56175 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13302 56176 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13303 5529 5610 5506 VDDHV pch_18 l=0.44u w=1.3u
m13304 5529 5854 56175 VDDHV pch_18 l=0.65u w=1.3u
m13305 5529 5854 56176 VDDHV pch_18 l=0.65u w=1.3u
m13306 5506 5610 5529 VDDHV pch_18 l=0.44u w=1.3u
m13307 5529 5610 5506 VDDHV pch_18 l=0.44u w=1.3u
m13308 56779 5854 5529 VDDHV pch_18 l=0.65u w=1.3u
m13309 56780 5854 5529 VDDHV pch_18 l=0.65u w=1.3u
m13310 5506 5610 5529 VDDHV pch_18 l=0.44u w=1.3u
m13311 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13312 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13313 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13314 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13315 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13316 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13317 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13318 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13319 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13320 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13321 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13322 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13323 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13324 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13325 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13326 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13327 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13328 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13329 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13330 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13331 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13332 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13333 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13334 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13335 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13336 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13337 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13338 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13339 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13340 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13341 VDDHV 5854 56779 VDDHV pch_18 l=0.65u w=1.3u
m13342 VDDHV 5854 56780 VDDHV pch_18 l=0.65u w=1.3u
m13343 57560 5610 5610 VDDHV pch_18 l=0.65u w=1.3u
m13344 57561 5610 5610 VDDHV pch_18 l=0.65u w=1.3u
m13345 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13346 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13347 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13348 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13349 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13350 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13351 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13352 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13353 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13354 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13355 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13356 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13357 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13358 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13359 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13360 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13361 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13362 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13363 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13364 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13365 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13366 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13367 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13368 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13369 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13370 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13371 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13372 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13373 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13374 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13375 5659 5610 57560 VDDHV pch_18 l=0.65u w=1.3u
m13376 5659 5610 57561 VDDHV pch_18 l=0.65u w=1.3u
m13377 58128 5610 5659 VDDHV pch_18 l=0.65u w=1.3u
m13378 58129 5610 5659 VDDHV pch_18 l=0.65u w=1.3u
m13379 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13380 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13381 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13382 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13383 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13384 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13385 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13386 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13387 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13388 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13389 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13390 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13391 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13392 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13393 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13394 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13395 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13396 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13397 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13398 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13399 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13400 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13401 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13402 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13403 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13404 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13405 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13406 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13407 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13408 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13409 VDDHV 5610 58128 VDDHV pch_18 l=0.65u w=1.3u
m13410 VDDHV 5610 58129 VDDHV pch_18 l=0.65u w=1.3u
m13411 58944 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13412 58945 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13413 5733 5610 5726 VDDHV pch_18 l=0.44u w=1.3u
m13414 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13415 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13416 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13417 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13418 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13419 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13420 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13421 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13422 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13423 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13424 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13425 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13426 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13427 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13428 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13429 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13430 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13431 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13432 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13433 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13434 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13435 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13436 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13437 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13438 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13439 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13440 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13441 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13442 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13443 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13444 5733 5854 58944 VDDHV pch_18 l=0.65u w=1.3u
m13445 5733 5854 58945 VDDHV pch_18 l=0.65u w=1.3u
m13446 5726 5610 5733 VDDHV pch_18 l=0.44u w=1.3u
m13447 5733 5610 5726 VDDHV pch_18 l=0.44u w=1.3u
m13448 59493 5854 5733 VDDHV pch_18 l=0.65u w=1.3u
m13449 59494 5854 5733 VDDHV pch_18 l=0.65u w=1.3u
m13450 5726 5610 5733 VDDHV pch_18 l=0.44u w=1.3u
m13451 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13452 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13453 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13454 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13455 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13456 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13457 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13458 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13459 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13460 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13461 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13462 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13463 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13464 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13465 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13466 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13467 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13468 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13469 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13470 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13471 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13472 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13473 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13474 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13475 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13476 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13477 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13478 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13479 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13480 VDDHV 4861 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13481 VDDHV 5854 59493 VDDHV pch_18 l=0.65u w=1.3u
m13482 VDDHV 5854 59494 VDDHV pch_18 l=0.65u w=1.3u
m13483 60605 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13484 60606 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13485 5139 5854 60605 VDDHV pch_18 l=0.65u w=1.3u
m13486 5139 5854 60606 VDDHV pch_18 l=0.65u w=1.3u
m13487 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13488 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13489 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13490 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13491 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13492 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13493 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13494 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13495 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13496 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13497 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13498 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13499 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13500 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13501 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13502 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13503 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13504 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13505 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13506 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13507 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13508 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13509 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13510 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13511 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13512 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13513 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13514 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13515 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13516 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13517 61446 5854 5139 VDDHV pch_18 l=0.65u w=1.3u
m13518 61447 5854 5139 VDDHV pch_18 l=0.65u w=1.3u
m13519 VDDHV 5854 61446 VDDHV pch_18 l=0.65u w=1.3u
m13520 VDDHV 5854 61447 VDDHV pch_18 l=0.65u w=1.3u
m13521 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13522 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13523 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13524 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13525 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13526 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13527 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13528 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13529 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13530 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13531 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13532 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13533 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13534 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13535 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13536 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13537 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13538 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13539 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13540 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13541 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13542 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13543 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13544 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13545 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13546 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13547 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13548 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13549 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13550 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13551 62465 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13552 62466 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13553 5040 5854 62465 VDDHV pch_18 l=0.65u w=1.3u
m13554 5040 5854 62466 VDDHV pch_18 l=0.65u w=1.3u
m13555 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13556 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13557 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13558 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13559 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13560 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13561 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13562 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13563 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13564 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13565 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13566 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13567 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13568 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13569 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13570 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13571 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13572 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13573 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13574 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13575 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13576 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13577 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13578 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13579 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13580 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13581 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13582 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13583 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13584 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13585 63430 5854 5040 VDDHV pch_18 l=0.65u w=1.3u
m13586 63431 5854 5040 VDDHV pch_18 l=0.65u w=1.3u
m13587 VDDHV 5854 63430 VDDHV pch_18 l=0.65u w=1.3u
m13588 VDDHV 5854 63431 VDDHV pch_18 l=0.65u w=1.3u
m13589 VDDHV 5643 5643 VDDHV pch_18 l=0.65u w=0.975u
m13590 5830 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13591 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13592 5645 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13593 VDDHV 2 5615 VDDHV pch_18 l=0.65u w=0.975u
m13594 5442 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13595 VDDHV 2 5411 VDDHV pch_18 l=0.65u w=0.975u
m13596 5412 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13597 VDDHV 2 5443 VDDHV pch_18 l=0.65u w=0.975u
m13598 5616 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13599 VDDHV 2 5646 VDDHV pch_18 l=0.65u w=0.975u
m13600 5816 5786 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13601 VDDHV 5786 5816 VDDHV pch_18 l=0.65u w=0.975u
m13602 5803 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13603 VDDHV 5643 5643 VDDHV pch_18 l=0.65u w=0.975u
m13604 5804 5067 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13605 VDDHV 5067 5804 VDDHV pch_18 l=0.65u w=0.975u
m13606 5647 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13607 VDDHV 2 5617 VDDHV pch_18 l=0.65u w=0.975u
m13608 5444 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13609 VDDHV 2 5413 VDDHV pch_18 l=0.65u w=0.975u
m13610 5414 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13611 VDDHV 2 5445 VDDHV pch_18 l=0.65u w=0.975u
m13612 5618 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13613 VDDHV 2 5648 VDDHV pch_18 l=0.65u w=0.975u
m13614 5774 5067 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13615 VDDHV 5067 5774 VDDHV pch_18 l=0.65u w=0.975u
m13616 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13617 VDDHV 5643 5643 VDDHV pch_18 l=0.65u w=0.975u
m13618 5775 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13619 VDDHV 2 5775 VDDHV pch_18 l=0.65u w=0.975u
m13620 5649 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13621 VDDHV 2 5619 VDDHV pch_18 l=0.65u w=0.975u
m13622 5446 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13623 VDDHV 2 5415 VDDHV pch_18 l=0.65u w=0.975u
m13624 5416 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13625 VDDHV 2 5447 VDDHV pch_18 l=0.65u w=0.975u
m13626 5620 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13627 VDDHV 2 5650 VDDHV pch_18 l=0.65u w=0.975u
m13628 5776 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13629 VDDHV 2 5776 VDDHV pch_18 l=0.65u w=0.975u
m13630 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13631 VDDHV 5643 5643 VDDHV pch_18 l=0.65u w=0.975u
m13632 5777 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13633 VDDHV 2 5777 VDDHV pch_18 l=0.65u w=0.975u
m13634 5651 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13635 VDDHV 2 5621 VDDHV pch_18 l=0.65u w=0.975u
m13636 5448 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13637 VDDHV 2 5417 VDDHV pch_18 l=0.65u w=0.975u
m13638 5418 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13639 VDDHV 2 5449 VDDHV pch_18 l=0.65u w=0.975u
m13640 5622 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13641 VDDHV 2 5652 VDDHV pch_18 l=0.65u w=0.975u
m13642 5778 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13643 VDDHV 2 5778 VDDHV pch_18 l=0.65u w=0.975u
m13644 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13645 VDDHV 5643 5643 VDDHV pch_18 l=0.65u w=0.975u
m13646 5779 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13647 VDDHV 2 5779 VDDHV pch_18 l=0.65u w=0.975u
m13648 5653 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13649 VDDHV 2 5623 VDDHV pch_18 l=0.65u w=0.975u
m13650 5450 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13651 VDDHV 2 5419 VDDHV pch_18 l=0.65u w=0.975u
m13652 5420 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13653 VDDHV 2 5451 VDDHV pch_18 l=0.65u w=0.975u
m13654 5624 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13655 VDDHV 2 5654 VDDHV pch_18 l=0.65u w=0.975u
m13656 5780 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13657 VDDHV 2 5780 VDDHV pch_18 l=0.65u w=0.975u
m13658 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13659 VDDHV 5643 5643 VDDHV pch_18 l=0.65u w=0.975u
m13660 5781 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13661 VDDHV 2 5781 VDDHV pch_18 l=0.65u w=0.975u
m13662 5655 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13663 VDDHV 2 5625 VDDHV pch_18 l=0.65u w=0.975u
m13664 5452 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13665 VDDHV 2 5421 VDDHV pch_18 l=0.65u w=0.975u
m13666 5422 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13667 VDDHV 2 5453 VDDHV pch_18 l=0.65u w=0.975u
m13668 5626 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13669 VDDHV 2 5656 VDDHV pch_18 l=0.65u w=0.975u
m13670 5782 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13671 VDDHV 2 5782 VDDHV pch_18 l=0.65u w=0.975u
m13672 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13673 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13674 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13675 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13676 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13677 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13678 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13679 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13680 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13681 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13682 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13683 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13684 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13685 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13686 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13687 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13688 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13689 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13690 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13691 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13692 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13693 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13694 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13695 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13696 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13697 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13698 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13699 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13700 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13701 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13702 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13703 63911 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13704 63912 5854 VDDHV VDDHV pch_18 l=0.65u w=1.3u
m13705 5860 5610 5854 VDDHV pch_18 l=0.44u w=1.3u
m13706 5860 5854 63911 VDDHV pch_18 l=0.65u w=1.3u
m13707 5860 5854 63912 VDDHV pch_18 l=0.65u w=1.3u
m13708 5854 5610 5860 VDDHV pch_18 l=0.44u w=1.3u
m13709 VDDHV 2 5815 VDDHV pch_18 l=0.65u w=0.975u
m13710 5858 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13711 VDDHV 2 5753 VDDHV pch_18 l=0.65u w=0.975u
m13712 5677 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13713 VDDHV 2 5582 VDDHV pch_18 l=0.65u w=0.975u
m13714 5474 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13715 VDDHV 2 5380 VDDHV pch_18 l=0.65u w=0.975u
m13716 5381 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13717 VDDHV 2 5475 VDDHV pch_18 l=0.65u w=0.975u
m13718 5583 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13719 VDDHV 2 5678 VDDHV pch_18 l=0.65u w=0.975u
m13720 5754 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13721 VDDHV 2 5595 VDDHV pch_18 l=0.65u w=0.975u
m13722 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13723 VDDHV 2 5595 VDDHV pch_18 l=0.65u w=0.975u
m13724 5804 5067 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13725 VDDHV 2 5755 VDDHV pch_18 l=0.65u w=0.975u
m13726 5679 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13727 VDDHV 2 5584 VDDHV pch_18 l=0.65u w=0.975u
m13728 5476 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13729 VDDHV 2 5382 VDDHV pch_18 l=0.65u w=0.975u
m13730 5383 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13731 VDDHV 2 5477 VDDHV pch_18 l=0.65u w=0.975u
m13732 5585 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13733 VDDHV 2 5680 VDDHV pch_18 l=0.65u w=0.975u
m13734 5756 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13735 VDDHV 5067 5774 VDDHV pch_18 l=0.65u w=0.975u
m13736 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13737 VDDHV 2 5595 VDDHV pch_18 l=0.65u w=0.975u
m13738 5775 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13739 VDDHV 2 5757 VDDHV pch_18 l=0.65u w=0.975u
m13740 5681 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13741 VDDHV 2 5586 VDDHV pch_18 l=0.65u w=0.975u
m13742 5478 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13743 VDDHV 2 5384 VDDHV pch_18 l=0.65u w=0.975u
m13744 5385 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13745 VDDHV 2 5479 VDDHV pch_18 l=0.65u w=0.975u
m13746 5587 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13747 VDDHV 2 5682 VDDHV pch_18 l=0.65u w=0.975u
m13748 5758 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13749 VDDHV 2 5776 VDDHV pch_18 l=0.65u w=0.975u
m13750 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13751 VDDHV 2 5595 VDDHV pch_18 l=0.65u w=0.975u
m13752 5777 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13753 VDDHV 2 5759 VDDHV pch_18 l=0.65u w=0.975u
m13754 5683 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13755 VDDHV 2 5588 VDDHV pch_18 l=0.65u w=0.975u
m13756 5480 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13757 VDDHV 2 5386 VDDHV pch_18 l=0.65u w=0.975u
m13758 5387 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13759 VDDHV 2 5481 VDDHV pch_18 l=0.65u w=0.975u
m13760 5589 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13761 VDDHV 2 5684 VDDHV pch_18 l=0.65u w=0.975u
m13762 5760 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13763 VDDHV 2 5778 VDDHV pch_18 l=0.65u w=0.975u
m13764 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13765 VDDHV 2 5595 VDDHV pch_18 l=0.65u w=0.975u
m13766 5779 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13767 VDDHV 2 5761 VDDHV pch_18 l=0.65u w=0.975u
m13768 5685 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13769 VDDHV 2 5590 VDDHV pch_18 l=0.65u w=0.975u
m13770 5482 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13771 VDDHV 2 5388 VDDHV pch_18 l=0.65u w=0.975u
m13772 5389 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13773 VDDHV 2 5483 VDDHV pch_18 l=0.65u w=0.975u
m13774 5591 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13775 VDDHV 2 5686 VDDHV pch_18 l=0.65u w=0.975u
m13776 5762 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13777 VDDHV 2 5780 VDDHV pch_18 l=0.65u w=0.975u
m13778 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13779 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13780 5781 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13781 VDDHV 2 5763 VDDHV pch_18 l=0.65u w=0.975u
m13782 5687 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13783 VDDHV 2 5592 VDDHV pch_18 l=0.65u w=0.975u
m13784 5484 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13785 VDDHV 2 5390 VDDHV pch_18 l=0.65u w=0.975u
m13786 5391 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13787 VDDHV 2 5485 VDDHV pch_18 l=0.65u w=0.975u
m13788 5593 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13789 VDDHV 2 5688 VDDHV pch_18 l=0.65u w=0.975u
m13790 5764 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13791 VDDHV 2 5782 VDDHV pch_18 l=0.65u w=0.975u
m13792 VDDHV 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13793 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13794 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13795 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13796 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13797 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13798 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13799 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13800 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13801 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13802 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13803 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13804 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13805 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13806 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13807 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13808 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13809 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13810 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13811 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13812 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13813 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13814 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13815 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13816 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13817 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13818 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13819 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13820 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13821 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13822 VDDHV 2 VDDHV VDDHV pch_18 l=1.9u w=2.98u
m13823 5860 5610 5854 VDDHV pch_18 l=0.44u w=1.3u
m13824 64199 5854 5860 VDDHV pch_18 l=0.65u w=1.3u
m13825 64200 5854 5860 VDDHV pch_18 l=0.65u w=1.3u
m13826 5854 5610 5860 VDDHV pch_18 l=0.44u w=1.3u
m13827 VDDHV 5854 64199 VDDHV pch_18 l=0.65u w=1.3u
m13828 VDDHV 5854 64200 VDDHV pch_18 l=0.65u w=1.3u
m13829 VDDHV 2 5814 VDDHV pch_18 l=0.65u w=0.975u
m13830 5823 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13831 VDDHV 2 5734 VDDHV pch_18 l=0.65u w=0.975u
m13832 5709 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13833 VDDHV 2 5551 VDDHV pch_18 l=0.65u w=0.975u
m13834 5513 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13835 VDDHV 2 5344 VDDHV pch_18 l=0.65u w=0.975u
m13836 5345 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13837 VDDHV 2 5514 VDDHV pch_18 l=0.65u w=0.975u
m13838 5552 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13839 VDDHV 2 5710 VDDHV pch_18 l=0.65u w=0.975u
m13840 5735 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13841 VDDHV 2 5595 VDDHV pch_18 l=0.65u w=0.975u
m13842 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13843 VDDHV 2 5595 VDDHV pch_18 l=0.65u w=0.975u
m13844 5595 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13845 VDDHV 2 5736 VDDHV pch_18 l=0.65u w=0.975u
m13846 5711 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13847 VDDHV 2 5553 VDDHV pch_18 l=0.65u w=0.975u
m13848 5515 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13849 VDDHV 2 5346 VDDHV pch_18 l=0.65u w=0.975u
m13850 5347 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13851 VDDHV 2 5516 VDDHV pch_18 l=0.65u w=0.975u
m13852 5554 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13853 VDDHV 2 5712 VDDHV pch_18 l=0.65u w=0.975u
m13854 5737 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13855 VDDHV 5067 5774 VDDHV pch_18 l=0.65u w=0.975u
m13856 5774 5067 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13857 VDDHV 2 5775 VDDHV pch_18 l=0.65u w=0.975u
m13858 5775 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13859 VDDHV 2 5738 VDDHV pch_18 l=0.65u w=0.975u
m13860 5713 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13861 VDDHV 2 5555 VDDHV pch_18 l=0.65u w=0.975u
m13862 5517 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13863 VDDHV 2 5348 VDDHV pch_18 l=0.65u w=0.975u
m13864 5349 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13865 VDDHV 2 5518 VDDHV pch_18 l=0.65u w=0.975u
m13866 5556 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13867 VDDHV 2 5714 VDDHV pch_18 l=0.65u w=0.975u
m13868 5739 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13869 VDDHV 2 5776 VDDHV pch_18 l=0.65u w=0.975u
m13870 5776 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13871 VDDHV 2 5777 VDDHV pch_18 l=0.65u w=0.975u
m13872 5777 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13873 VDDHV 2 5740 VDDHV pch_18 l=0.65u w=0.975u
m13874 5715 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13875 VDDHV 2 5557 VDDHV pch_18 l=0.65u w=0.975u
m13876 5519 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13877 VDDHV 2 5350 VDDHV pch_18 l=0.65u w=0.975u
m13878 5351 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13879 VDDHV 2 5520 VDDHV pch_18 l=0.65u w=0.975u
m13880 5558 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13881 VDDHV 2 5716 VDDHV pch_18 l=0.65u w=0.975u
m13882 5741 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13883 VDDHV 2 5778 VDDHV pch_18 l=0.65u w=0.975u
m13884 5778 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13885 VDDHV 2 5779 VDDHV pch_18 l=0.65u w=0.975u
m13886 5779 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13887 VDDHV 2 5742 VDDHV pch_18 l=0.65u w=0.975u
m13888 5717 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13889 VDDHV 2 5559 VDDHV pch_18 l=0.65u w=0.975u
m13890 5521 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13891 VDDHV 2 5352 VDDHV pch_18 l=0.65u w=0.975u
m13892 5353 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13893 VDDHV 2 5522 VDDHV pch_18 l=0.65u w=0.975u
m13894 5560 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13895 VDDHV 2 5718 VDDHV pch_18 l=0.65u w=0.975u
m13896 5743 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13897 VDDHV 2 5780 VDDHV pch_18 l=0.65u w=0.975u
m13898 5780 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13899 VDDHV 2 5781 VDDHV pch_18 l=0.65u w=0.975u
m13900 5781 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13901 VDDHV 2 5744 VDDHV pch_18 l=0.65u w=0.975u
m13902 5719 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13903 VDDHV 2 5561 VDDHV pch_18 l=0.65u w=0.975u
m13904 5523 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13905 VDDHV 2 5354 VDDHV pch_18 l=0.65u w=0.975u
m13906 5355 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13907 VDDHV 2 5524 VDDHV pch_18 l=0.65u w=0.975u
m13908 5562 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13909 VDDHV 2 5720 VDDHV pch_18 l=0.65u w=0.975u
m13910 5745 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13911 VDDHV 2 5782 VDDHV pch_18 l=0.65u w=0.975u
m13912 5782 2 VDDHV VDDHV pch_18 l=0.65u w=0.975u
m13913 6 PD VDDREF VDDREF pch l=0.04u w=0.8u
m13914 9 6 VDDREF VDDREF pch l=0.04u w=0.12u
m13915 VDDREF FREF 9 VDDREF pch l=0.04u w=0.4u
m13916 9 FREF VDDREF VDDREF pch l=0.04u w=0.4u
m13917 10 FREF VDDREF VDDREF pch l=0.04u w=0.8u
m13918 11 9 VDDREF VDDREF pch l=0.04u w=0.8u
m13919 12 10 VDDREF VDDREF pch l=0.04u w=0.8u
m13920 VDDREF 9 11 VDDREF pch l=0.04u w=0.8u
m13921 VDDREF 10 12 VDDREF pch l=0.04u w=0.8u
m13922 11 9 VDDREF VDDREF pch l=0.04u w=0.8u
m13923 12 10 VDDREF VDDREF pch l=0.04u w=0.8u
m13924 VDDREF 9 11 VDDREF pch l=0.04u w=0.8u
m13925 VDDREF 10 12 VDDREF pch l=0.04u w=0.8u
m13926 27284 REFDIV[3] VDDREF VDDREF pch l=0.04u w=0.8u
m13927 16 212 VDDREF VDDREF pch l=0.04u w=0.8u
m13928 VDDREF 30 14 VDDREF pch l=0.04u w=0.8u
m13929 17 110 VDDREF VDDREF pch l=0.04u w=0.8u
m13930 18 66 VDDREF VDDREF pch l=0.04u w=0.8u
m13931 27309 REFDIV[4] 27284 VDDREF pch l=0.04u w=0.8u
m13932 VDDREF 11 16 VDDREF pch l=0.04u w=0.8u
m13933 VDDREF 91 17 VDDREF pch l=0.04u w=0.8u
m13934 VDDREF 94 18 VDDREF pch l=0.04u w=0.8u
m13935 15 REFDIV[5] 27309 VDDREF pch l=0.04u w=0.8u
m13936 16 11 VDDREF VDDREF pch l=0.04u w=0.8u
m13937 VDDREF 19 20 VDDREF pch l=0.04u w=1u
m13938 35 138 VDDREF VDDREF pch l=0.04u w=0.8u
m13939 21 77 VDDREF VDDREF pch l=0.04u w=0.8u
m13940 36 130 VDDREF VDDREF pch l=0.04u w=0.8u
m13941 37 139 VDDREF VDDREF pch l=0.04u w=0.8u
m13942 22 78 VDDREF VDDREF pch l=0.04u w=0.8u
m13943 38 140 VDDREF VDDREF pch l=0.04u w=0.8u
m13944 39 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m13945 40 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m13946 VDDREF 23 24 VDDREF pch l=0.04u w=1u
m13947 41 141 VDDREF VDDREF pch l=0.04u w=0.8u
m13948 25 79 VDDREF VDDREF pch l=0.04u w=0.8u
m13949 42 FRAC[0] VDDREF VDDREF pch l=0.04u w=0.8u
m13950 43 60 VDDREF VDDREF pch l=0.04u w=0.8u
m13951 44 61 VDDREF VDDREF pch l=0.04u w=0.8u
m13952 VDDREF 109 26 VDDREF pch l=0.04u w=0.8u
m13953 27 81 VDDREF VDDREF pch l=0.04u w=0.8u
m13954 45 132 VDDREF VDDREF pch l=0.04u w=0.8u
m13955 46 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m13956 47 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m13957 48 145 VDDREF VDDREF pch l=0.04u w=0.8u
m13958 28 82 VDDREF VDDREF pch l=0.04u w=0.8u
m13959 49 146 VDDREF VDDREF pch l=0.04u w=0.8u
m13960 50 26 VDDREF VDDREF pch l=0.04u w=0.8u
m13961 51 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m13962 52 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m13963 53 141 VDDREF VDDREF pch l=0.04u w=0.8u
m13964 29 83 VDDREF VDDREF pch l=0.04u w=0.8u
m13965 54 FRAC[0] VDDREF VDDREF pch l=0.04u w=0.8u
m13966 55 26 VDDREF VDDREF pch l=0.04u w=0.8u
m13967 30 84 VDDREF VDDREF pch l=0.04u w=0.8u
m13968 VDDREF 31 32 VDDREF pch l=0.04u w=1u
m13969 VDDREF 34 33 VDDREF pch l=0.04u w=1u
m13970 VDDREF 125 35 VDDREF pch l=0.04u w=0.8u
m13971 VDDREF 246 21 VDDREF pch l=0.04u w=0.8u
m13972 VDDREF 126 36 VDDREF pch l=0.04u w=0.8u
m13973 VDDREF 127 37 VDDREF pch l=0.04u w=0.8u
m13974 VDDREF 247 22 VDDREF pch l=0.04u w=0.8u
m13975 VDDREF 128 38 VDDREF pch l=0.04u w=0.8u
m13976 VDDREF 298 39 VDDREF pch l=0.04u w=0.8u
m13977 VDDREF 299 40 VDDREF pch l=0.04u w=0.8u
m13978 VDDREF 129 41 VDDREF pch l=0.04u w=0.8u
m13979 VDDREF 248 25 VDDREF pch l=0.04u w=0.8u
m13980 VDDREF 130 42 VDDREF pch l=0.04u w=0.8u
m13981 VDDREF 249 27 VDDREF pch l=0.04u w=0.8u
m13982 VDDREF 131 45 VDDREF pch l=0.04u w=0.8u
m13983 VDDREF 132 48 VDDREF pch l=0.04u w=0.8u
m13984 VDDREF 250 28 VDDREF pch l=0.04u w=0.8u
m13985 VDDREF 133 49 VDDREF pch l=0.04u w=0.8u
m13986 VDDREF 134 50 VDDREF pch l=0.04u w=0.8u
m13987 VDDREF 135 53 VDDREF pch l=0.04u w=0.8u
m13988 VDDREF 251 29 VDDREF pch l=0.04u w=0.8u
m13989 VDDREF 136 54 VDDREF pch l=0.04u w=0.8u
m13990 VDDREF FBDIV[0] 55 VDDREF pch l=0.04u w=0.8u
m13991 VDDREF 2648 30 VDDREF pch l=0.04u w=0.8u
m13992 VDDREF 56 57 VDDREF pch l=0.04u w=1u
m13993 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m13994 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m13995 67 91 VDDREF VDDREF pch l=0.04u w=0.8u
m13996 68 94 VDDREF VDDREF pch l=0.04u w=0.8u
m13997 27358 REFDIV[1] VDDREF VDDREF pch l=0.04u w=0.8u
m13998 76 16 VDDREF VDDREF pch l=0.04u w=0.8u
m13999 58 69 60 VDDREF pch l=0.04u w=0.8u
m14000 59 70 61 VDDREF pch l=0.04u w=0.8u
m14001 80 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14002 71 4328 62 VDDREF pch l=0.04u w=0.8u
m14003 72 4328 63 VDDREF pch l=0.04u w=0.8u
m14004 73 4328 64 VDDREF pch l=0.04u w=0.8u
m14005 74 4328 65 VDDREF pch l=0.04u w=0.8u
m14006 VDDREF 110 66 VDDREF pch l=0.04u w=0.8u
m14007 VDDREF 231 VDDREF VDDREF pch l=0.26u w=1u
m14008 VDDREF 234 VDDREF VDDREF pch l=0.26u w=1u
m14009 75 REFDIV[2] 27358 VDDREF pch l=0.04u w=0.8u
m14010 VDDREF 16 76 VDDREF pch l=0.04u w=0.8u
m14011 92 125 VDDREF VDDREF pch l=0.04u w=0.8u
m14012 VDDREF 1159 77 VDDREF pch l=0.04u w=0.8u
m14013 93 126 VDDREF VDDREF pch l=0.04u w=0.8u
m14014 95 127 VDDREF VDDREF pch l=0.04u w=0.8u
m14015 VDDREF 1162 78 VDDREF pch l=0.04u w=0.8u
m14016 96 128 VDDREF VDDREF pch l=0.04u w=0.8u
m14017 97 39 VDDREF VDDREF pch l=0.04u w=0.8u
m14018 98 40 VDDREF VDDREF pch l=0.04u w=0.8u
m14019 99 129 VDDREF VDDREF pch l=0.04u w=0.8u
m14020 VDDREF 1165 79 VDDREF pch l=0.04u w=0.8u
m14021 100 130 VDDREF VDDREF pch l=0.04u w=0.8u
m14022 69 60 58 VDDREF pch l=0.04u w=0.8u
m14023 70 61 59 VDDREF pch l=0.04u w=0.8u
m14024 VDDREF 131 81 VDDREF pch l=0.04u w=0.8u
m14025 101 131 VDDREF VDDREF pch l=0.04u w=0.8u
m14026 27367 46 71 VDDREF pch l=0.04u w=0.12u
m14027 27368 47 72 VDDREF pch l=0.04u w=0.12u
m14028 102 132 VDDREF VDDREF pch l=0.04u w=0.8u
m14029 VDDREF 1169 82 VDDREF pch l=0.04u w=0.8u
m14030 103 133 VDDREF VDDREF pch l=0.04u w=0.8u
m14031 104 134 VDDREF VDDREF pch l=0.04u w=0.8u
m14032 27369 51 73 VDDREF pch l=0.04u w=0.12u
m14033 27370 52 74 VDDREF pch l=0.04u w=0.12u
m14034 105 135 VDDREF VDDREF pch l=0.04u w=0.8u
m14035 VDDREF 1173 83 VDDREF pch l=0.04u w=0.8u
m14036 106 136 VDDREF VDDREF pch l=0.04u w=0.8u
m14037 107 FBDIV[0] VDDREF VDDREF pch l=0.04u w=0.8u
m14038 VDDREF 154 84 VDDREF pch l=0.04u w=0.8u
m14039 108 DSMPD VDDREF VDDREF pch l=0.04u w=0.8u
m14040 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14041 VDDREF 86 85 VDDREF pch l=0.04u w=1u
m14042 VDDREF 87 88 VDDREF pch l=0.04u w=1u
m14043 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m14044 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m14045 76 16 VDDREF VDDREF pch l=0.04u w=0.8u
m14046 89 110 91 VDDREF pch l=0.04u w=0.8u
m14047 77 311 VDDREF VDDREF pch l=0.04u w=0.8u
m14048 90 66 94 VDDREF pch l=0.04u w=0.8u
m14049 78 312 VDDREF VDDREF pch l=0.04u w=0.8u
m14050 79 314 VDDREF VDDREF pch l=0.04u w=0.8u
m14051 81 316 VDDREF VDDREF pch l=0.04u w=0.8u
m14052 VDDREF 143 27367 VDDREF pch l=0.04u w=0.12u
m14053 VDDREF 144 27368 VDDREF pch l=0.04u w=0.12u
m14054 82 317 VDDREF VDDREF pch l=0.04u w=0.8u
m14055 VDDREF 147 27369 VDDREF pch l=0.04u w=0.12u
m14056 VDDREF 148 27370 VDDREF pch l=0.04u w=0.12u
m14057 83 319 VDDREF VDDREF pch l=0.04u w=0.8u
m14058 27387 14 VDDREF VDDREF pch l=0.04u w=0.24u
m14059 117 4328 109 VDDREF pch l=0.04u w=0.8u
m14060 VDDREF 231 VDDREF VDDREF pch l=0.26u w=1u
m14061 VDDREF 234 VDDREF VDDREF pch l=0.26u w=1u
m14062 VDDREF 16 76 VDDREF pch l=0.04u w=0.8u
m14063 110 91 89 VDDREF pch l=0.04u w=0.8u
m14064 VDDREF 160 77 VDDREF pch l=0.04u w=0.8u
m14065 66 94 90 VDDREF pch l=0.04u w=0.8u
m14066 VDDREF 162 78 VDDREF pch l=0.04u w=0.8u
m14067 VDDREF 163 79 VDDREF pch l=0.04u w=0.8u
m14068 VDDREF 164 81 VDDREF pch l=0.04u w=0.8u
m14069 143 71 VDDREF VDDREF pch l=0.04u w=0.8u
m14070 144 72 VDDREF VDDREF pch l=0.04u w=0.8u
m14071 VDDREF 165 82 VDDREF pch l=0.04u w=0.8u
m14072 147 73 VDDREF VDDREF pch l=0.04u w=0.8u
m14073 148 74 VDDREF VDDREF pch l=0.04u w=0.8u
m14074 VDDREF 166 83 VDDREF pch l=0.04u w=0.8u
m14075 149 75 VDDREF VDDREF pch l=0.04u w=0.8u
m14076 154 886 27387 VDDREF pch l=0.04u w=0.24u
m14077 150 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14078 151 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14079 111 138 125 VDDREF pch l=0.04u w=0.8u
m14080 112 130 126 VDDREF pch l=0.04u w=0.8u
m14081 113 139 127 VDDREF pch l=0.04u w=0.8u
m14082 114 140 128 VDDREF pch l=0.04u w=0.8u
m14083 152 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14084 153 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14085 115 141 129 VDDREF pch l=0.04u w=0.8u
m14086 116 FRAC[0] 130 VDDREF pch l=0.04u w=0.8u
m14087 27398 80 117 VDDREF pch l=0.04u w=0.12u
m14088 118 132 131 VDDREF pch l=0.04u w=0.8u
m14089 119 145 132 VDDREF pch l=0.04u w=0.8u
m14090 120 146 133 VDDREF pch l=0.04u w=0.8u
m14091 121 26 134 VDDREF pch l=0.04u w=0.8u
m14092 122 141 135 VDDREF pch l=0.04u w=0.8u
m14093 123 FRAC[0] 136 VDDREF pch l=0.04u w=0.8u
m14094 124 26 FBDIV[0] VDDREF pch l=0.04u w=0.8u
m14095 155 14 VDDREF VDDREF pch l=0.04u w=0.8u
m14096 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14097 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14098 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14099 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m14100 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m14101 156 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14102 157 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14103 76 16 VDDREF VDDREF pch l=0.04u w=0.8u
m14104 VDDREF 15 149 VDDREF pch l=0.04u w=0.8u
m14105 158 270 154 VDDREF pch l=0.04u w=0.8u
m14106 138 125 111 VDDREF pch l=0.04u w=0.8u
m14107 130 126 112 VDDREF pch l=0.04u w=0.8u
m14108 139 127 113 VDDREF pch l=0.04u w=0.8u
m14109 140 128 114 VDDREF pch l=0.04u w=0.8u
m14110 141 129 115 VDDREF pch l=0.04u w=0.8u
m14111 FRAC[0] 130 116 VDDREF pch l=0.04u w=0.8u
m14112 VDDREF 177 27398 VDDREF pch l=0.04u w=0.12u
m14113 132 131 118 VDDREF pch l=0.04u w=0.8u
m14114 145 132 119 VDDREF pch l=0.04u w=0.8u
m14115 146 133 120 VDDREF pch l=0.04u w=0.8u
m14116 26 134 121 VDDREF pch l=0.04u w=0.8u
m14117 141 135 122 VDDREF pch l=0.04u w=0.8u
m14118 FRAC[0] 136 123 VDDREF pch l=0.04u w=0.8u
m14119 26 FBDIV[0] 124 VDDREF pch l=0.04u w=0.8u
m14120 VDDREF 108 155 VDDREF pch l=0.04u w=0.8u
m14121 VDDREF 231 VDDREF VDDREF pch l=0.26u w=1u
m14122 VDDREF 234 VDDREF VDDREF pch l=0.26u w=1u
m14123 VDDREF 16 76 VDDREF pch l=0.04u w=0.8u
m14124 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14125 159 89 VDDREF VDDREF pch l=0.04u w=0.8u
m14126 VDDREF 194 160 VDDREF pch l=0.04u w=0.8u
m14127 161 90 VDDREF VDDREF pch l=0.04u w=0.8u
m14128 VDDREF 195 162 VDDREF pch l=0.04u w=0.8u
m14129 VDDREF 196 163 VDDREF pch l=0.04u w=0.8u
m14130 177 117 VDDREF VDDREF pch l=0.04u w=0.8u
m14131 VDDREF 197 164 VDDREF pch l=0.04u w=0.8u
m14132 169 46 143 VDDREF pch l=0.04u w=0.8u
m14133 170 47 144 VDDREF pch l=0.04u w=0.8u
m14134 VDDREF 198 165 VDDREF pch l=0.04u w=0.8u
m14135 171 51 147 VDDREF pch l=0.04u w=0.8u
m14136 172 52 148 VDDREF pch l=0.04u w=0.8u
m14137 VDDREF 199 166 VDDREF pch l=0.04u w=0.8u
m14138 173 4328 167 VDDREF pch l=0.04u w=0.8u
m14139 174 4328 168 VDDREF pch l=0.04u w=0.8u
m14140 175 4328 97 VDDREF pch l=0.04u w=0.8u
m14141 176 4328 98 VDDREF pch l=0.04u w=0.8u
m14142 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14143 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14144 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m14145 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m14146 76 16 VDDREF VDDREF pch l=0.04u w=0.8u
m14147 191 4328 58 VDDREF pch l=0.04u w=0.8u
m14148 192 4328 59 VDDREF pch l=0.04u w=0.8u
m14149 VDDREF 110 159 VDDREF pch l=0.04u w=0.8u
m14150 VDDREF 293 161 VDDREF pch l=0.04u w=0.8u
m14151 27423 4328 169 VDDREF pch l=0.04u w=0.12u
m14152 27424 4328 170 VDDREF pch l=0.04u w=0.12u
m14153 27425 4328 171 VDDREF pch l=0.04u w=0.12u
m14154 27426 4328 172 VDDREF pch l=0.04u w=0.12u
m14155 193 149 VDDREF VDDREF pch l=0.04u w=0.8u
m14156 158 217 VDDREF VDDREF pch l=0.04u w=0.8u
m14157 27427 150 173 VDDREF pch l=0.04u w=0.12u
m14158 27428 151 174 VDDREF pch l=0.04u w=0.12u
m14159 178 111 VDDREF VDDREF pch l=0.04u w=0.8u
m14160 179 112 VDDREF VDDREF pch l=0.04u w=0.8u
m14161 180 113 VDDREF VDDREF pch l=0.04u w=0.8u
m14162 181 114 VDDREF VDDREF pch l=0.04u w=0.8u
m14163 27429 152 175 VDDREF pch l=0.04u w=0.12u
m14164 27430 153 176 VDDREF pch l=0.04u w=0.12u
m14165 182 115 VDDREF VDDREF pch l=0.04u w=0.8u
m14166 183 116 VDDREF VDDREF pch l=0.04u w=0.8u
m14167 184 118 VDDREF VDDREF pch l=0.04u w=0.8u
m14168 185 119 VDDREF VDDREF pch l=0.04u w=0.8u
m14169 186 120 VDDREF VDDREF pch l=0.04u w=0.8u
m14170 187 121 VDDREF VDDREF pch l=0.04u w=0.8u
m14171 188 122 VDDREF VDDREF pch l=0.04u w=0.8u
m14172 189 123 VDDREF VDDREF pch l=0.04u w=0.8u
m14173 190 124 VDDREF VDDREF pch l=0.04u w=0.8u
m14174 200 155 VDDREF VDDREF pch l=0.04u w=0.8u
m14175 VDDREF 231 VDDREF VDDREF pch l=0.26u w=1u
m14176 VDDREF 234 VDDREF VDDREF pch l=0.26u w=1u
m14177 VDDREF 16 76 VDDREF pch l=0.04u w=0.8u
m14178 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14179 27434 156 191 VDDREF pch l=0.04u w=0.12u
m14180 27435 157 192 VDDREF pch l=0.04u w=0.12u
m14181 VDDREF 202 27423 VDDREF pch l=0.04u w=0.12u
m14182 VDDREF 203 27424 VDDREF pch l=0.04u w=0.12u
m14183 VDDREF 204 27425 VDDREF pch l=0.04u w=0.12u
m14184 VDDREF 205 27426 VDDREF pch l=0.04u w=0.12u
m14185 VDDREF 2648 158 VDDREF pch l=0.04u w=0.8u
m14186 VDDREF 207 27427 VDDREF pch l=0.04u w=0.12u
m14187 VDDREF 208 27428 VDDREF pch l=0.04u w=0.12u
m14188 VDDREF 21 178 VDDREF pch l=0.04u w=0.8u
m14189 VDDREF 610 194 VDDREF pch l=0.04u w=0.8u
m14190 VDDREF 110 179 VDDREF pch l=0.04u w=0.8u
m14191 VDDREF 22 180 VDDREF pch l=0.04u w=0.8u
m14192 VDDREF 611 195 VDDREF pch l=0.04u w=0.8u
m14193 VDDREF 313 181 VDDREF pch l=0.04u w=0.8u
m14194 VDDREF 210 27429 VDDREF pch l=0.04u w=0.12u
m14195 VDDREF 211 27430 VDDREF pch l=0.04u w=0.12u
m14196 VDDREF 25 182 VDDREF pch l=0.04u w=0.8u
m14197 VDDREF 612 196 VDDREF pch l=0.04u w=0.8u
m14198 VDDREF 315 183 VDDREF pch l=0.04u w=0.8u
m14199 201 80 177 VDDREF pch l=0.04u w=0.8u
m14200 VDDREF 613 197 VDDREF pch l=0.04u w=0.8u
m14201 VDDREF 27 184 VDDREF pch l=0.04u w=0.8u
m14202 VDDREF 28 185 VDDREF pch l=0.04u w=0.8u
m14203 VDDREF 614 198 VDDREF pch l=0.04u w=0.8u
m14204 VDDREF 131 186 VDDREF pch l=0.04u w=0.8u
m14205 VDDREF 318 187 VDDREF pch l=0.04u w=0.8u
m14206 VDDREF 29 188 VDDREF pch l=0.04u w=0.8u
m14207 VDDREF 615 199 VDDREF pch l=0.04u w=0.8u
m14208 VDDREF 131 189 VDDREF pch l=0.04u w=0.8u
m14209 VDDREF 318 190 VDDREF pch l=0.04u w=0.8u
m14210 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14211 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14212 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m14213 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m14214 VDDREF 214 27434 VDDREF pch l=0.04u w=0.12u
m14215 VDDREF 215 27435 VDDREF pch l=0.04u w=0.12u
m14216 202 169 VDDREF VDDREF pch l=0.04u w=0.8u
m14217 203 170 VDDREF VDDREF pch l=0.04u w=0.8u
m14218 204 171 VDDREF VDDREF pch l=0.04u w=0.8u
m14219 205 172 VDDREF VDDREF pch l=0.04u w=0.8u
m14220 27447 158 VDDREF VDDREF pch l=0.04u w=0.12u
m14221 206 159 VDDREF VDDREF pch l=0.04u w=0.8u
m14222 207 173 VDDREF VDDREF pch l=0.04u w=0.8u
m14223 208 174 VDDREF VDDREF pch l=0.04u w=0.8u
m14224 194 903 VDDREF VDDREF pch l=0.04u w=0.8u
m14225 209 161 VDDREF VDDREF pch l=0.04u w=0.8u
m14226 195 904 VDDREF VDDREF pch l=0.04u w=0.8u
m14227 210 175 VDDREF VDDREF pch l=0.04u w=0.8u
m14228 211 176 VDDREF VDDREF pch l=0.04u w=0.8u
m14229 196 905 VDDREF VDDREF pch l=0.04u w=0.8u
m14230 27448 4328 201 VDDREF pch l=0.04u w=0.12u
m14231 197 906 VDDREF VDDREF pch l=0.04u w=0.8u
m14232 198 907 VDDREF VDDREF pch l=0.04u w=0.8u
m14233 199 908 VDDREF VDDREF pch l=0.04u w=0.8u
m14234 27449 PD VDDREF VDDREF pch l=0.04u w=0.8u
m14235 VDDREF 231 VDDREF VDDREF pch l=0.26u w=1u
m14236 VDDREF 234 VDDREF VDDREF pch l=0.26u w=1u
m14237 213 155 VDDREF VDDREF pch l=0.04u w=0.8u
m14238 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14239 214 191 VDDREF VDDREF pch l=0.04u w=0.8u
m14240 215 192 VDDREF VDDREF pch l=0.04u w=0.8u
m14241 216 236 VDDREF VDDREF pch l=0.04u w=0.8u
m14242 217 270 27447 VDDREF pch l=0.04u w=0.12u
m14243 VDDREF 17 206 VDDREF pch l=0.04u w=0.8u
m14244 VDDREF 1190 194 VDDREF pch l=0.04u w=0.8u
m14245 VDDREF 18 209 VDDREF pch l=0.04u w=0.8u
m14246 VDDREF 1191 195 VDDREF pch l=0.04u w=0.8u
m14247 VDDREF 1192 196 VDDREF pch l=0.04u w=0.8u
m14248 VDDREF 241 27448 VDDREF pch l=0.04u w=0.12u
m14249 VDDREF 1193 197 VDDREF pch l=0.04u w=0.8u
m14250 VDDREF 1194 198 VDDREF pch l=0.04u w=0.8u
m14251 VDDREF 1195 199 VDDREF pch l=0.04u w=0.8u
m14252 212 193 27449 VDDREF pch l=0.04u w=0.8u
m14253 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14254 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14255 218 178 VDDREF VDDREF pch l=0.04u w=0.8u
m14256 219 179 VDDREF VDDREF pch l=0.04u w=0.8u
m14257 220 180 VDDREF VDDREF pch l=0.04u w=0.8u
m14258 221 181 VDDREF VDDREF pch l=0.04u w=0.8u
m14259 222 182 VDDREF VDDREF pch l=0.04u w=0.8u
m14260 223 183 VDDREF VDDREF pch l=0.04u w=0.8u
m14261 224 184 VDDREF VDDREF pch l=0.04u w=0.8u
m14262 225 185 VDDREF VDDREF pch l=0.04u w=0.8u
m14263 226 186 VDDREF VDDREF pch l=0.04u w=0.8u
m14264 227 187 VDDREF VDDREF pch l=0.04u w=0.8u
m14265 228 188 VDDREF VDDREF pch l=0.04u w=0.8u
m14266 229 189 VDDREF VDDREF pch l=0.04u w=0.8u
m14267 230 190 VDDREF VDDREF pch l=0.04u w=0.8u
m14268 232 232 VDDREF VDDREF pch l=0.04u w=1u
m14269 233 233 VDDREF VDDREF pch l=0.04u w=1u
m14270 VDDREF FBDIV[0] 213 VDDREF pch l=0.04u w=0.8u
m14271 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m14272 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m14273 235 259 216 VDDREF pch l=0.04u w=0.8u
m14274 VDDREF 886 217 VDDREF pch l=0.04u w=0.8u
m14275 241 201 VDDREF VDDREF pch l=0.04u w=0.8u
m14276 242 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14277 243 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14278 244 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14279 245 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14280 237 150 207 VDDREF pch l=0.04u w=0.8u
m14281 238 151 208 VDDREF pch l=0.04u w=0.8u
m14282 VDDREF 35 218 VDDREF pch l=0.04u w=0.8u
m14283 VDDREF 36 219 VDDREF pch l=0.04u w=0.8u
m14284 VDDREF 37 220 VDDREF pch l=0.04u w=0.8u
m14285 VDDREF 38 221 VDDREF pch l=0.04u w=0.8u
m14286 239 152 210 VDDREF pch l=0.04u w=0.8u
m14287 240 153 211 VDDREF pch l=0.04u w=0.8u
m14288 VDDREF 41 222 VDDREF pch l=0.04u w=0.8u
m14289 VDDREF 42 223 VDDREF pch l=0.04u w=0.8u
m14290 VDDREF 45 224 VDDREF pch l=0.04u w=0.8u
m14291 VDDREF 48 225 VDDREF pch l=0.04u w=0.8u
m14292 VDDREF 49 226 VDDREF pch l=0.04u w=0.8u
m14293 VDDREF 50 227 VDDREF pch l=0.04u w=0.8u
m14294 VDDREF 53 228 VDDREF pch l=0.04u w=0.8u
m14295 VDDREF 54 229 VDDREF pch l=0.04u w=0.8u
m14296 VDDREF 55 230 VDDREF pch l=0.04u w=0.8u
m14297 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14298 259 216 235 VDDREF pch l=0.04u w=0.8u
m14299 257 156 214 VDDREF pch l=0.04u w=0.8u
m14300 258 157 215 VDDREF pch l=0.04u w=0.8u
m14301 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14302 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14303 260 89 VDDREF VDDREF pch l=0.04u w=0.8u
m14304 27468 4328 237 VDDREF pch l=0.04u w=0.12u
m14305 27469 4328 238 VDDREF pch l=0.04u w=0.12u
m14306 VDDREF 353 246 VDDREF pch l=0.04u w=0.8u
m14307 261 90 VDDREF VDDREF pch l=0.04u w=0.8u
m14308 VDDREF 356 247 VDDREF pch l=0.04u w=0.8u
m14309 27470 4328 239 VDDREF pch l=0.04u w=0.12u
m14310 27471 4328 240 VDDREF pch l=0.04u w=0.12u
m14311 VDDREF 361 248 VDDREF pch l=0.04u w=0.8u
m14312 VDDREF 363 249 VDDREF pch l=0.04u w=0.8u
m14313 VDDREF 366 250 VDDREF pch l=0.04u w=0.8u
m14314 VDDREF 370 251 VDDREF pch l=0.04u w=0.8u
m14315 236 212 VDDREF VDDREF pch l=0.04u w=0.8u
m14316 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m14317 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m14318 VDDREF 252 253 VDDREF pch l=0.04u w=1u
m14319 VDDREF 255 254 VDDREF pch l=0.04u w=1u
m14320 265 200 VDDREF VDDREF pch l=0.04u w=0.8u
m14321 27476 4328 257 VDDREF pch l=0.04u w=0.12u
m14322 27477 4328 258 VDDREF pch l=0.04u w=0.12u
m14323 270 886 VDDREF VDDREF pch l=0.04u w=0.8u
m14324 VDDREF 292 27468 VDDREF pch l=0.04u w=0.12u
m14325 VDDREF 126 27469 VDDREF pch l=0.04u w=0.12u
m14326 VDDREF 294 27470 VDDREF pch l=0.04u w=0.12u
m14327 VDDREF 130 27471 VDDREF pch l=0.04u w=0.12u
m14328 266 4328 262 VDDREF pch l=0.04u w=0.8u
m14329 267 4328 263 VDDREF pch l=0.04u w=0.8u
m14330 268 4328 264 VDDREF pch l=0.04u w=0.8u
m14331 269 4328 134 VDDREF pch l=0.04u w=0.8u
m14332 273 111 VDDREF VDDREF pch l=0.04u w=0.8u
m14333 275 112 VDDREF VDDREF pch l=0.04u w=0.8u
m14334 276 113 VDDREF VDDREF pch l=0.04u w=0.8u
m14335 278 114 VDDREF VDDREF pch l=0.04u w=0.8u
m14336 279 115 VDDREF VDDREF pch l=0.04u w=0.8u
m14337 281 116 VDDREF VDDREF pch l=0.04u w=0.8u
m14338 283 118 VDDREF VDDREF pch l=0.04u w=0.8u
m14339 284 119 VDDREF VDDREF pch l=0.04u w=0.8u
m14340 286 120 VDDREF VDDREF pch l=0.04u w=0.8u
m14341 287 121 VDDREF VDDREF pch l=0.04u w=0.8u
m14342 288 122 VDDREF VDDREF pch l=0.04u w=0.8u
m14343 290 123 VDDREF VDDREF pch l=0.04u w=0.8u
m14344 291 124 VDDREF VDDREF pch l=0.04u w=0.8u
m14345 VDDREF 241 265 VDDREF pch l=0.04u w=0.8u
m14346 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14347 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14348 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14349 VDDREF 304 27476 VDDREF pch l=0.04u w=0.12u
m14350 VDDREF 305 27477 VDDREF pch l=0.04u w=0.12u
m14351 292 237 VDDREF VDDREF pch l=0.04u w=0.8u
m14352 126 238 VDDREF VDDREF pch l=0.04u w=0.8u
m14353 VDDREF 307 VDDREF VDDREF pch l=0.26u w=1u
m14354 294 239 VDDREF VDDREF pch l=0.04u w=0.8u
m14355 130 240 VDDREF VDDREF pch l=0.04u w=0.8u
m14356 VDDREF 309 VDDREF VDDREF pch l=0.26u w=1u
m14357 27484 242 266 VDDREF pch l=0.04u w=0.12u
m14358 27485 243 267 VDDREF pch l=0.04u w=0.12u
m14359 27486 244 268 VDDREF pch l=0.04u w=0.12u
m14360 27487 245 269 VDDREF pch l=0.04u w=0.12u
m14361 VDDREF 447 VDDREF VDDREF pch l=0.26u w=1u
m14362 VDDREF 450 VDDREF VDDREF pch l=0.26u w=1u
m14363 271 110 89 VDDREF pch l=0.04u w=0.8u
m14364 167 311 274 VDDREF pch l=0.04u w=0.8u
m14365 272 293 90 VDDREF pch l=0.04u w=0.8u
m14366 298 312 277 VDDREF pch l=0.04u w=0.8u
m14367 300 314 280 VDDREF pch l=0.04u w=0.8u
m14368 301 316 282 VDDREF pch l=0.04u w=0.8u
m14369 63 317 285 VDDREF pch l=0.04u w=0.8u
m14370 65 319 289 VDDREF pch l=0.04u w=0.8u
m14371 303 485 VDDREF VDDREF pch l=0.04u w=0.8u
m14372 304 257 VDDREF VDDREF pch l=0.04u w=0.8u
m14373 305 258 VDDREF VDDREF pch l=0.04u w=0.8u
m14374 306 377 VDDREF VDDREF pch l=0.04u w=0.8u
m14375 308 308 VDDREF VDDREF pch l=0.04u w=1u
m14376 310 310 VDDREF VDDREF pch l=0.04u w=1u
m14377 VDDREF 323 27484 VDDREF pch l=0.04u w=0.12u
m14378 VDDREF 324 27485 VDDREF pch l=0.04u w=0.12u
m14379 VDDREF 325 27486 VDDREF pch l=0.04u w=0.12u
m14380 VDDREF 326 27487 VDDREF pch l=0.04u w=0.12u
m14381 VDDREF 327 LOCK VDDREF pch l=0.04u w=0.8u
m14382 110 89 271 VDDREF pch l=0.04u w=0.8u
m14383 311 274 167 VDDREF pch l=0.04u w=0.8u
m14384 293 90 272 VDDREF pch l=0.04u w=0.8u
m14385 312 277 298 VDDREF pch l=0.04u w=0.8u
m14386 314 280 300 VDDREF pch l=0.04u w=0.8u
m14387 316 282 301 VDDREF pch l=0.04u w=0.8u
m14388 317 285 63 VDDREF pch l=0.04u w=0.8u
m14389 319 289 65 VDDREF pch l=0.04u w=0.8u
m14390 VDDREF 485 303 VDDREF pch l=0.04u w=0.8u
m14391 296 21 111 VDDREF pch l=0.04u w=0.8u
m14392 168 110 112 VDDREF pch l=0.04u w=0.8u
m14393 297 22 113 VDDREF pch l=0.04u w=0.8u
m14394 299 313 114 VDDREF pch l=0.04u w=0.8u
m14395 127 25 115 VDDREF pch l=0.04u w=0.8u
m14396 128 315 116 VDDREF pch l=0.04u w=0.8u
m14397 109 27 118 VDDREF pch l=0.04u w=0.8u
m14398 263 28 119 VDDREF pch l=0.04u w=0.8u
m14399 302 131 120 VDDREF pch l=0.04u w=0.8u
m14400 145 318 121 VDDREF pch l=0.04u w=0.8u
m14401 134 29 122 VDDREF pch l=0.04u w=0.8u
m14402 146 131 123 VDDREF pch l=0.04u w=0.8u
m14403 141 318 124 VDDREF pch l=0.04u w=0.8u
m14404 320 265 VDDREF VDDREF pch l=0.04u w=0.8u
m14405 VDDREF 334 VDDREF VDDREF pch l=0.26u w=1u
m14406 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14407 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14408 VDDREF 447 VDDREF VDDREF pch l=0.26u w=1u
m14409 VDDREF 450 VDDREF VDDREF pch l=0.26u w=1u
m14410 323 266 VDDREF VDDREF pch l=0.04u w=0.8u
m14411 324 267 VDDREF VDDREF pch l=0.04u w=0.8u
m14412 325 268 VDDREF VDDREF pch l=0.04u w=0.8u
m14413 326 269 VDDREF VDDREF pch l=0.04u w=0.8u
m14414 303 485 VDDREF VDDREF pch l=0.04u w=0.8u
m14415 21 111 296 VDDREF pch l=0.04u w=0.8u
m14416 110 112 168 VDDREF pch l=0.04u w=0.8u
m14417 22 113 297 VDDREF pch l=0.04u w=0.8u
m14418 313 114 299 VDDREF pch l=0.04u w=0.8u
m14419 25 115 127 VDDREF pch l=0.04u w=0.8u
m14420 315 116 128 VDDREF pch l=0.04u w=0.8u
m14421 27 118 109 VDDREF pch l=0.04u w=0.8u
m14422 28 119 263 VDDREF pch l=0.04u w=0.8u
m14423 131 120 302 VDDREF pch l=0.04u w=0.8u
m14424 318 121 145 VDDREF pch l=0.04u w=0.8u
m14425 29 122 134 VDDREF pch l=0.04u w=0.8u
m14426 131 123 146 VDDREF pch l=0.04u w=0.8u
m14427 318 124 141 VDDREF pch l=0.04u w=0.8u
m14428 VDDREF 213 320 VDDREF pch l=0.04u w=0.8u
m14429 335 335 VDDREF VDDREF pch l=0.04u w=1u
m14430 VDDREF 304 321 VDDREF pch l=0.04u w=0.8u
m14431 VDDREF 305 322 VDDREF pch l=0.04u w=0.8u
m14432 336 377 VDDREF VDDREF pch l=0.04u w=0.8u
m14433 VDDREF 485 303 VDDREF pch l=0.04u w=0.8u
m14434 327 378 VDDREF VDDREF pch l=0.04u w=0.8u
m14435 337 415 VDDREF VDDREF pch l=0.04u w=0.8u
m14436 VDDREF 311 328 VDDREF pch l=0.04u w=0.8u
m14437 338 379 VDDREF VDDREF pch l=0.04u w=0.8u
m14438 VDDREF 312 329 VDDREF pch l=0.04u w=0.8u
m14439 VDDREF 314 330 VDDREF pch l=0.04u w=0.8u
m14440 VDDREF 316 331 VDDREF pch l=0.04u w=0.8u
m14441 VDDREF 317 332 VDDREF pch l=0.04u w=0.8u
m14442 VDDREF 319 333 VDDREF pch l=0.04u w=0.8u
m14443 VDDREF 374 VDDREF VDDREF pch l=0.26u w=1u
m14444 VDDREF 375 VDDREF VDDREF pch l=0.26u w=1u
m14445 VDDREF 447 VDDREF VDDREF pch l=0.26u w=1u
m14446 VDDREF 450 VDDREF VDDREF pch l=0.26u w=1u
m14447 346 321 VDDREF VDDREF pch l=0.04u w=0.8u
m14448 347 322 VDDREF VDDREF pch l=0.04u w=0.8u
m14449 VDDREF REFDIV[0] 336 VDDREF pch l=0.04u w=0.8u
m14450 348 242 323 VDDREF pch l=0.04u w=0.8u
m14451 349 243 324 VDDREF pch l=0.04u w=0.8u
m14452 350 244 325 VDDREF pch l=0.04u w=0.8u
m14453 351 245 326 VDDREF pch l=0.04u w=0.8u
m14454 VDDREF 2648 327 VDDREF pch l=0.04u w=0.8u
m14455 VDDREF 395 337 VDDREF pch l=0.04u w=0.8u
m14456 VDDREF 398 338 VDDREF pch l=0.04u w=0.8u
m14457 VDDREF 339 340 VDDREF pch l=0.04u w=1u
m14458 352 458 VDDREF VDDREF pch l=0.04u w=0.8u
m14459 354 442 VDDREF VDDREF pch l=0.04u w=0.8u
m14460 355 139 VDDREF VDDREF pch l=0.04u w=0.8u
m14461 357 459 VDDREF VDDREF pch l=0.04u w=0.8u
m14462 358 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m14463 359 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m14464 VDDREF 341 342 VDDREF pch l=0.04u w=1u
m14465 360 460 VDDREF VDDREF pch l=0.04u w=0.8u
m14466 362 FRAC[1] VDDREF VDDREF pch l=0.04u w=0.8u
m14467 VDDREF 412 343 VDDREF pch l=0.04u w=0.8u
m14468 364 443 VDDREF VDDREF pch l=0.04u w=0.8u
m14469 365 462 VDDREF VDDREF pch l=0.04u w=0.8u
m14470 367 264 VDDREF VDDREF pch l=0.04u w=0.8u
m14471 368 343 VDDREF VDDREF pch l=0.04u w=0.8u
m14472 369 460 VDDREF VDDREF pch l=0.04u w=0.8u
m14473 371 FRAC[1] VDDREF VDDREF pch l=0.04u w=0.8u
m14474 372 343 VDDREF VDDREF pch l=0.04u w=0.8u
m14475 VDDREF 344 345 VDDREF pch l=0.04u w=1u
m14476 373 373 VDDREF VDDREF pch l=0.04u w=1u
m14477 376 376 VDDREF VDDREF pch l=0.04u w=1u
m14478 27526 4328 348 VDDREF pch l=0.04u w=0.12u
m14479 27527 4328 349 VDDREF pch l=0.04u w=0.12u
m14480 27528 4328 350 VDDREF pch l=0.04u w=0.12u
m14481 27529 4328 351 VDDREF pch l=0.04u w=0.12u
m14482 377 457 VDDREF VDDREF pch l=0.04u w=0.8u
m14483 VDDREF 437 352 VDDREF pch l=0.04u w=0.8u
m14484 353 530 VDDREF VDDREF pch l=0.04u w=0.8u
m14485 VDDREF 438 354 VDDREF pch l=0.04u w=0.8u
m14486 VDDREF 439 355 VDDREF pch l=0.04u w=0.8u
m14487 356 533 VDDREF VDDREF pch l=0.04u w=0.8u
m14488 VDDREF 440 357 VDDREF pch l=0.04u w=0.8u
m14489 VDDREF 597 358 VDDREF pch l=0.04u w=0.8u
m14490 VDDREF 598 359 VDDREF pch l=0.04u w=0.8u
m14491 VDDREF 441 360 VDDREF pch l=0.04u w=0.8u
m14492 361 536 VDDREF VDDREF pch l=0.04u w=0.8u
m14493 VDDREF 442 362 VDDREF pch l=0.04u w=0.8u
m14494 363 538 VDDREF VDDREF pch l=0.04u w=0.8u
m14495 VDDREF 131 364 VDDREF pch l=0.04u w=0.8u
m14496 VDDREF 443 365 VDDREF pch l=0.04u w=0.8u
m14497 366 541 VDDREF VDDREF pch l=0.04u w=0.8u
m14498 VDDREF 391 367 VDDREF pch l=0.04u w=0.8u
m14499 VDDREF 444 368 VDDREF pch l=0.04u w=0.8u
m14500 VDDREF 445 369 VDDREF pch l=0.04u w=0.8u
m14501 370 545 VDDREF VDDREF pch l=0.04u w=0.8u
m14502 VDDREF 392 371 VDDREF pch l=0.04u w=0.8u
m14503 VDDREF FBDIV[1] 372 VDDREF pch l=0.04u w=0.8u
m14504 VDDREF 447 VDDREF VDDREF pch l=0.26u w=1u
m14505 VDDREF 450 VDDREF VDDREF pch l=0.26u w=1u
m14506 385 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14507 386 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14508 VDDREF 391 27526 VDDREF pch l=0.04u w=0.12u
m14509 VDDREF 132 27527 VDDREF pch l=0.04u w=0.12u
m14510 VDDREF 392 27528 VDDREF pch l=0.04u w=0.12u
m14511 VDDREF 135 27529 VDDREF pch l=0.04u w=0.12u
m14512 387 306 VDDREF VDDREF pch l=0.04u w=0.8u
m14513 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14514 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14515 VDDREF 457 377 VDDREF pch l=0.04u w=0.8u
m14516 VDDREF 416 378 VDDREF pch l=0.04u w=0.8u
m14517 388 395 VDDREF VDDREF pch l=0.04u w=0.8u
m14518 VDDREF 418 353 VDDREF pch l=0.04u w=0.8u
m14519 389 398 VDDREF VDDREF pch l=0.04u w=0.8u
m14520 VDDREF 421 356 VDDREF pch l=0.04u w=0.8u
m14521 VDDREF 424 361 VDDREF pch l=0.04u w=0.8u
m14522 VDDREF 427 363 VDDREF pch l=0.04u w=0.8u
m14523 VDDREF 430 366 VDDREF pch l=0.04u w=0.8u
m14524 VDDREF 434 370 VDDREF pch l=0.04u w=0.8u
m14525 390 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14526 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14527 VDDREF 1918 379 VDDREF pch l=0.04u w=0.8u
m14528 VDDREF 381 380 VDDREF pch l=0.04u w=1u
m14529 VDDREF 382 383 VDDREF pch l=0.04u w=1u
m14530 391 348 VDDREF VDDREF pch l=0.04u w=0.8u
m14531 132 349 VDDREF VDDREF pch l=0.04u w=0.8u
m14532 392 350 VDDREF VDDREF pch l=0.04u w=0.8u
m14533 135 351 VDDREF VDDREF pch l=0.04u w=0.8u
m14534 VDDREF 235 387 VDDREF pch l=0.04u w=0.8u
m14535 377 457 VDDREF VDDREF pch l=0.04u w=0.8u
m14536 27546 LOCK VDDREF VDDREF pch l=0.04u w=0.24u
m14537 396 437 VDDREF VDDREF pch l=0.04u w=0.8u
m14538 397 438 VDDREF VDDREF pch l=0.04u w=0.8u
m14539 399 439 VDDREF VDDREF pch l=0.04u w=0.8u
m14540 400 440 VDDREF VDDREF pch l=0.04u w=0.8u
m14541 401 358 VDDREF VDDREF pch l=0.04u w=0.8u
m14542 402 359 VDDREF VDDREF pch l=0.04u w=0.8u
m14543 403 441 VDDREF VDDREF pch l=0.04u w=0.8u
m14544 404 442 VDDREF VDDREF pch l=0.04u w=0.8u
m14545 405 131 VDDREF VDDREF pch l=0.04u w=0.8u
m14546 406 443 VDDREF VDDREF pch l=0.04u w=0.8u
m14547 407 391 VDDREF VDDREF pch l=0.04u w=0.8u
m14548 408 444 VDDREF VDDREF pch l=0.04u w=0.8u
m14549 409 445 VDDREF VDDREF pch l=0.04u w=0.8u
m14550 410 392 VDDREF VDDREF pch l=0.04u w=0.8u
m14551 411 FBDIV[1] VDDREF VDDREF pch l=0.04u w=0.8u
m14552 VDDREF 447 VDDREF VDDREF pch l=0.26u w=1u
m14553 VDDREF 450 VDDREF VDDREF pch l=0.26u w=1u
m14554 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14555 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14556 413 4328 304 VDDREF pch l=0.04u w=0.8u
m14557 414 4328 305 VDDREF pch l=0.04u w=0.8u
m14558 VDDREF 457 377 VDDREF pch l=0.04u w=0.8u
m14559 416 605 27546 VDDREF pch l=0.04u w=0.24u
m14560 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14561 393 415 395 VDDREF pch l=0.04u w=0.8u
m14562 418 274 VDDREF VDDREF pch l=0.04u w=0.8u
m14563 394 379 398 VDDREF pch l=0.04u w=0.8u
m14564 421 277 VDDREF VDDREF pch l=0.04u w=0.8u
m14565 424 280 VDDREF VDDREF pch l=0.04u w=0.8u
m14566 427 282 VDDREF VDDREF pch l=0.04u w=0.8u
m14567 430 285 VDDREF VDDREF pch l=0.04u w=0.8u
m14568 434 289 VDDREF VDDREF pch l=0.04u w=0.8u
m14569 426 4328 412 VDDREF pch l=0.04u w=0.8u
m14570 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14571 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14572 448 448 VDDREF VDDREF pch l=0.04u w=1u
m14573 449 449 VDDREF VDDREF pch l=0.04u w=1u
m14574 27559 385 413 VDDREF pch l=0.04u w=0.12u
m14575 27560 386 414 VDDREF pch l=0.04u w=0.12u
m14576 451 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14577 452 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14578 453 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14579 454 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14580 455 387 VDDREF VDDREF pch l=0.04u w=0.8u
m14581 456 561 416 VDDREF pch l=0.04u w=0.8u
m14582 415 395 393 VDDREF pch l=0.04u w=0.8u
m14583 VDDREF 311 418 VDDREF pch l=0.04u w=0.8u
m14584 379 398 394 VDDREF pch l=0.04u w=0.8u
m14585 VDDREF 312 421 VDDREF pch l=0.04u w=0.8u
m14586 VDDREF 314 424 VDDREF pch l=0.04u w=0.8u
m14587 VDDREF 316 427 VDDREF pch l=0.04u w=0.8u
m14588 VDDREF 317 430 VDDREF pch l=0.04u w=0.8u
m14589 VDDREF 319 434 VDDREF pch l=0.04u w=0.8u
m14590 463 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14591 464 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14592 417 458 437 VDDREF pch l=0.04u w=0.8u
m14593 419 442 438 VDDREF pch l=0.04u w=0.8u
m14594 420 139 439 VDDREF pch l=0.04u w=0.8u
m14595 422 459 440 VDDREF pch l=0.04u w=0.8u
m14596 465 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14597 466 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14598 423 460 441 VDDREF pch l=0.04u w=0.8u
m14599 425 FRAC[1] 442 VDDREF pch l=0.04u w=0.8u
m14600 27561 390 426 VDDREF pch l=0.04u w=0.12u
m14601 428 443 131 VDDREF pch l=0.04u w=0.8u
m14602 429 462 443 VDDREF pch l=0.04u w=0.8u
m14603 431 264 391 VDDREF pch l=0.04u w=0.8u
m14604 432 343 444 VDDREF pch l=0.04u w=0.8u
m14605 433 460 445 VDDREF pch l=0.04u w=0.8u
m14606 435 FRAC[1] 392 VDDREF pch l=0.04u w=0.8u
m14607 436 343 FBDIV[1] VDDREF pch l=0.04u w=0.8u
m14608 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14609 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14610 VDDREF 479 27559 VDDREF pch l=0.04u w=0.12u
m14611 VDDREF 480 27560 VDDREF pch l=0.04u w=0.12u
m14612 VDDREF 336 455 VDDREF pch l=0.04u w=0.8u
m14613 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14614 VDDREF 508 457 VDDREF pch l=0.04u w=0.8u
m14615 458 437 417 VDDREF pch l=0.04u w=0.8u
m14616 442 438 419 VDDREF pch l=0.04u w=0.8u
m14617 139 439 420 VDDREF pch l=0.04u w=0.8u
m14618 459 440 422 VDDREF pch l=0.04u w=0.8u
m14619 460 441 423 VDDREF pch l=0.04u w=0.8u
m14620 FRAC[1] 442 425 VDDREF pch l=0.04u w=0.8u
m14621 VDDREF 490 27561 VDDREF pch l=0.04u w=0.12u
m14622 443 131 428 VDDREF pch l=0.04u w=0.8u
m14623 462 443 429 VDDREF pch l=0.04u w=0.8u
m14624 264 391 431 VDDREF pch l=0.04u w=0.8u
m14625 343 444 432 VDDREF pch l=0.04u w=0.8u
m14626 460 445 433 VDDREF pch l=0.04u w=0.8u
m14627 FRAC[1] 392 435 VDDREF pch l=0.04u w=0.8u
m14628 343 FBDIV[1] 436 VDDREF pch l=0.04u w=0.8u
m14629 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14630 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14631 VDDREF 467 468 VDDREF pch l=0.04u w=1u
m14632 VDDREF 470 469 VDDREF pch l=0.04u w=1u
m14633 479 413 VDDREF VDDREF pch l=0.04u w=0.8u
m14634 480 414 VDDREF VDDREF pch l=0.04u w=0.8u
m14635 455 336 VDDREF VDDREF pch l=0.04u w=0.8u
m14636 481 4328 471 VDDREF pch l=0.04u w=0.8u
m14637 482 4328 302 VDDREF pch l=0.04u w=0.8u
m14638 483 4328 472 VDDREF pch l=0.04u w=0.8u
m14639 484 4328 146 VDDREF pch l=0.04u w=0.8u
m14640 456 521 VDDREF VDDREF pch l=0.04u w=0.8u
m14641 473 393 VDDREF VDDREF pch l=0.04u w=0.8u
m14642 311 292 474 VDDREF pch l=0.04u w=0.8u
m14643 475 394 VDDREF VDDREF pch l=0.04u w=0.8u
m14644 312 300 139 VDDREF pch l=0.04u w=0.8u
m14645 314 294 FRAC[23] VDDREF pch l=0.04u w=0.8u
m14646 490 426 VDDREF VDDREF pch l=0.04u w=0.8u
m14647 316 347 203 VDDREF pch l=0.04u w=0.8u
m14648 317 203 65 VDDREF pch l=0.04u w=0.8u
m14649 319 205 FRAC[23] VDDREF pch l=0.04u w=0.8u
m14650 486 4328 477 VDDREF pch l=0.04u w=0.8u
m14651 487 4328 478 VDDREF pch l=0.04u w=0.8u
m14652 488 4328 401 VDDREF pch l=0.04u w=0.8u
m14653 489 4328 402 VDDREF pch l=0.04u w=0.8u
m14654 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14655 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14656 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14657 VDDREF 387 455 VDDREF pch l=0.04u w=0.8u
m14658 27579 451 481 VDDREF pch l=0.04u w=0.12u
m14659 27580 452 482 VDDREF pch l=0.04u w=0.12u
m14660 27581 453 483 VDDREF pch l=0.04u w=0.12u
m14661 27582 454 484 VDDREF pch l=0.04u w=0.12u
m14662 VDDREF 2648 456 VDDREF pch l=0.04u w=0.8u
m14663 VDDREF 508 485 VDDREF pch l=0.04u w=0.8u
m14664 VDDREF 206 473 VDDREF pch l=0.04u w=0.8u
m14665 292 474 311 VDDREF pch l=0.04u w=0.8u
m14666 VDDREF 209 475 VDDREF pch l=0.04u w=0.8u
m14667 300 139 312 VDDREF pch l=0.04u w=0.8u
m14668 294 FRAC[23] 314 VDDREF pch l=0.04u w=0.8u
m14669 347 203 316 VDDREF pch l=0.04u w=0.8u
m14670 203 65 317 VDDREF pch l=0.04u w=0.8u
m14671 205 FRAC[23] 319 VDDREF pch l=0.04u w=0.8u
m14672 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14673 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14674 27583 463 486 VDDREF pch l=0.04u w=0.12u
m14675 27584 464 487 VDDREF pch l=0.04u w=0.12u
m14676 491 417 VDDREF VDDREF pch l=0.04u w=0.8u
m14677 492 419 VDDREF VDDREF pch l=0.04u w=0.8u
m14678 493 420 VDDREF VDDREF pch l=0.04u w=0.8u
m14679 494 422 VDDREF VDDREF pch l=0.04u w=0.8u
m14680 27585 465 488 VDDREF pch l=0.04u w=0.12u
m14681 27586 466 489 VDDREF pch l=0.04u w=0.12u
m14682 495 423 VDDREF VDDREF pch l=0.04u w=0.8u
m14683 496 425 VDDREF VDDREF pch l=0.04u w=0.8u
m14684 497 428 VDDREF VDDREF pch l=0.04u w=0.8u
m14685 498 429 VDDREF VDDREF pch l=0.04u w=0.8u
m14686 499 431 VDDREF VDDREF pch l=0.04u w=0.8u
m14687 500 432 VDDREF VDDREF pch l=0.04u w=0.8u
m14688 501 433 VDDREF VDDREF pch l=0.04u w=0.8u
m14689 502 435 VDDREF VDDREF pch l=0.04u w=0.8u
m14690 503 436 VDDREF VDDREF pch l=0.04u w=0.8u
m14691 504 155 VDDREF VDDREF pch l=0.04u w=0.8u
m14692 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m14693 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m14694 505 385 479 VDDREF pch l=0.04u w=0.8u
m14695 506 386 480 VDDREF pch l=0.04u w=0.8u
m14696 VDDREF 516 27579 VDDREF pch l=0.04u w=0.12u
m14697 VDDREF 517 27580 VDDREF pch l=0.04u w=0.12u
m14698 VDDREF 518 27581 VDDREF pch l=0.04u w=0.12u
m14699 VDDREF 519 27582 VDDREF pch l=0.04u w=0.12u
m14700 27591 456 VDDREF VDDREF pch l=0.04u w=0.12u
m14701 VDDREF 523 27583 VDDREF pch l=0.04u w=0.12u
m14702 VDDREF 524 27584 VDDREF pch l=0.04u w=0.12u
m14703 VDDREF 218 491 VDDREF pch l=0.04u w=0.8u
m14704 VDDREF 219 492 VDDREF pch l=0.04u w=0.8u
m14705 VDDREF 220 493 VDDREF pch l=0.04u w=0.8u
m14706 VDDREF 221 494 VDDREF pch l=0.04u w=0.8u
m14707 VDDREF 526 27585 VDDREF pch l=0.04u w=0.12u
m14708 VDDREF 527 27586 VDDREF pch l=0.04u w=0.12u
m14709 VDDREF 222 495 VDDREF pch l=0.04u w=0.8u
m14710 VDDREF 223 496 VDDREF pch l=0.04u w=0.8u
m14711 507 390 490 VDDREF pch l=0.04u w=0.8u
m14712 VDDREF 224 497 VDDREF pch l=0.04u w=0.8u
m14713 VDDREF 225 498 VDDREF pch l=0.04u w=0.8u
m14714 VDDREF 226 499 VDDREF pch l=0.04u w=0.8u
m14715 VDDREF 227 500 VDDREF pch l=0.04u w=0.8u
m14716 VDDREF 228 501 VDDREF pch l=0.04u w=0.8u
m14717 VDDREF 229 502 VDDREF pch l=0.04u w=0.8u
m14718 VDDREF 230 503 VDDREF pch l=0.04u w=0.8u
m14719 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14720 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14721 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14722 27599 4328 505 VDDREF pch l=0.04u w=0.12u
m14723 27600 4328 506 VDDREF pch l=0.04u w=0.12u
m14724 516 481 VDDREF VDDREF pch l=0.04u w=0.8u
m14725 517 482 VDDREF VDDREF pch l=0.04u w=0.8u
m14726 518 483 VDDREF VDDREF pch l=0.04u w=0.8u
m14727 519 484 VDDREF VDDREF pch l=0.04u w=0.8u
m14728 520 76 VDDREF VDDREF pch l=0.04u w=0.8u
m14729 521 561 27591 VDDREF pch l=0.04u w=0.12u
m14730 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14731 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14732 508 560 VDDREF VDDREF pch l=0.04u w=0.8u
m14733 522 473 VDDREF VDDREF pch l=0.04u w=0.8u
m14734 523 486 VDDREF VDDREF pch l=0.04u w=0.8u
m14735 524 487 VDDREF VDDREF pch l=0.04u w=0.8u
m14736 VDDREF 292 509 VDDREF pch l=0.04u w=0.8u
m14737 525 475 VDDREF VDDREF pch l=0.04u w=0.8u
m14738 VDDREF 300 510 VDDREF pch l=0.04u w=0.8u
m14739 526 488 VDDREF VDDREF pch l=0.04u w=0.8u
m14740 527 489 VDDREF VDDREF pch l=0.04u w=0.8u
m14741 VDDREF 294 511 VDDREF pch l=0.04u w=0.8u
m14742 27602 4328 507 VDDREF pch l=0.04u w=0.12u
m14743 VDDREF 347 512 VDDREF pch l=0.04u w=0.8u
m14744 VDDREF 203 513 VDDREF pch l=0.04u w=0.8u
m14745 VDDREF 205 514 VDDREF pch l=0.04u w=0.8u
m14746 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m14747 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m14748 528 155 VDDREF VDDREF pch l=0.04u w=0.8u
m14749 VDDREF 548 27599 VDDREF pch l=0.04u w=0.12u
m14750 VDDREF 549 27600 VDDREF pch l=0.04u w=0.12u
m14751 VDDREF 605 521 VDDREF pch l=0.04u w=0.8u
m14752 VDDREF 764 508 VDDREF pch l=0.04u w=0.8u
m14753 VDDREF 337 522 VDDREF pch l=0.04u w=0.8u
m14754 VDDREF 338 525 VDDREF pch l=0.04u w=0.8u
m14755 VDDREF 559 27602 VDDREF pch l=0.04u w=0.12u
m14756 529 491 VDDREF VDDREF pch l=0.04u w=0.8u
m14757 531 492 VDDREF VDDREF pch l=0.04u w=0.8u
m14758 532 493 VDDREF VDDREF pch l=0.04u w=0.8u
m14759 534 494 VDDREF VDDREF pch l=0.04u w=0.8u
m14760 535 495 VDDREF VDDREF pch l=0.04u w=0.8u
m14761 537 496 VDDREF VDDREF pch l=0.04u w=0.8u
m14762 539 497 VDDREF VDDREF pch l=0.04u w=0.8u
m14763 540 498 VDDREF VDDREF pch l=0.04u w=0.8u
m14764 542 499 VDDREF VDDREF pch l=0.04u w=0.8u
m14765 543 500 VDDREF VDDREF pch l=0.04u w=0.8u
m14766 544 501 VDDREF VDDREF pch l=0.04u w=0.8u
m14767 546 502 VDDREF VDDREF pch l=0.04u w=0.8u
m14768 547 503 VDDREF VDDREF pch l=0.04u w=0.8u
m14769 VDDREF FBDIV[1] 528 VDDREF pch l=0.04u w=0.8u
m14770 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14771 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14772 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14773 548 505 VDDREF VDDREF pch l=0.04u w=0.8u
m14774 549 506 VDDREF VDDREF pch l=0.04u w=0.8u
m14775 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14776 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14777 550 451 516 VDDREF pch l=0.04u w=0.8u
m14778 551 452 517 VDDREF pch l=0.04u w=0.8u
m14779 552 453 518 VDDREF pch l=0.04u w=0.8u
m14780 553 454 519 VDDREF pch l=0.04u w=0.8u
m14781 554 76 455 VDDREF pch l=0.04u w=0.8u
m14782 559 507 VDDREF VDDREF pch l=0.04u w=0.8u
m14783 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m14784 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m14785 555 463 523 VDDREF pch l=0.04u w=0.8u
m14786 556 464 524 VDDREF pch l=0.04u w=0.8u
m14787 VDDREF 352 529 VDDREF pch l=0.04u w=0.8u
m14788 530 292 VDDREF VDDREF pch l=0.04u w=0.8u
m14789 VDDREF 354 531 VDDREF pch l=0.04u w=0.8u
m14790 VDDREF 355 532 VDDREF pch l=0.04u w=0.8u
m14791 533 300 VDDREF VDDREF pch l=0.04u w=0.8u
m14792 VDDREF 357 534 VDDREF pch l=0.04u w=0.8u
m14793 557 465 526 VDDREF pch l=0.04u w=0.8u
m14794 558 466 527 VDDREF pch l=0.04u w=0.8u
m14795 VDDREF 360 535 VDDREF pch l=0.04u w=0.8u
m14796 536 294 VDDREF VDDREF pch l=0.04u w=0.8u
m14797 VDDREF 362 537 VDDREF pch l=0.04u w=0.8u
m14798 538 347 VDDREF VDDREF pch l=0.04u w=0.8u
m14799 VDDREF 364 539 VDDREF pch l=0.04u w=0.8u
m14800 VDDREF 365 540 VDDREF pch l=0.04u w=0.8u
m14801 541 203 VDDREF VDDREF pch l=0.04u w=0.8u
m14802 VDDREF 367 542 VDDREF pch l=0.04u w=0.8u
m14803 VDDREF 368 543 VDDREF pch l=0.04u w=0.8u
m14804 VDDREF 369 544 VDDREF pch l=0.04u w=0.8u
m14805 545 205 VDDREF VDDREF pch l=0.04u w=0.8u
m14806 VDDREF 371 546 VDDREF pch l=0.04u w=0.8u
m14807 VDDREF 372 547 VDDREF pch l=0.04u w=0.8u
m14808 27615 4328 550 VDDREF pch l=0.04u w=0.12u
m14809 27616 4328 551 VDDREF pch l=0.04u w=0.12u
m14810 27617 4328 552 VDDREF pch l=0.04u w=0.12u
m14811 27618 4328 553 VDDREF pch l=0.04u w=0.12u
m14812 27620 520 554 VDDREF pch l=0.04u w=0.12u
m14813 561 605 VDDREF VDDREF pch l=0.04u w=0.8u
m14814 VDDREF 594 560 VDDREF pch l=0.04u w=0.8u
m14815 562 393 VDDREF VDDREF pch l=0.04u w=0.8u
m14816 27621 4328 555 VDDREF pch l=0.04u w=0.12u
m14817 27622 4328 556 VDDREF pch l=0.04u w=0.12u
m14818 VDDREF 474 530 VDDREF pch l=0.04u w=0.8u
m14819 563 394 VDDREF VDDREF pch l=0.04u w=0.8u
m14820 VDDREF 139 533 VDDREF pch l=0.04u w=0.8u
m14821 27623 4328 557 VDDREF pch l=0.04u w=0.12u
m14822 27624 4328 558 VDDREF pch l=0.04u w=0.12u
m14823 VDDREF FRAC[23] 536 VDDREF pch l=0.04u w=0.8u
m14824 VDDREF 203 538 VDDREF pch l=0.04u w=0.8u
m14825 VDDREF 65 541 VDDREF pch l=0.04u w=0.8u
m14826 VDDREF FRAC[23] 545 VDDREF pch l=0.04u w=0.8u
m14827 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14828 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14829 564 504 VDDREF VDDREF pch l=0.04u w=0.8u
m14830 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14831 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14832 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14833 565 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14834 566 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14835 VDDREF 589 27615 VDDREF pch l=0.04u w=0.12u
m14836 VDDREF 133 27616 VDDREF pch l=0.04u w=0.12u
m14837 VDDREF 590 27617 VDDREF pch l=0.04u w=0.12u
m14838 VDDREF 136 27618 VDDREF pch l=0.04u w=0.12u
m14839 VDDREF 591 27620 VDDREF pch l=0.04u w=0.12u
m14840 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m14841 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m14842 27633 485 VDDREF VDDREF pch l=0.04u w=0.24u
m14843 VDDREF 592 27621 VDDREF pch l=0.04u w=0.12u
m14844 VDDREF 438 27622 VDDREF pch l=0.04u w=0.12u
m14845 VDDREF 593 27623 VDDREF pch l=0.04u w=0.12u
m14846 VDDREF 442 27624 VDDREF pch l=0.04u w=0.12u
m14847 570 417 VDDREF VDDREF pch l=0.04u w=0.8u
m14848 572 419 VDDREF VDDREF pch l=0.04u w=0.8u
m14849 573 420 VDDREF VDDREF pch l=0.04u w=0.8u
m14850 575 422 VDDREF VDDREF pch l=0.04u w=0.8u
m14851 576 423 VDDREF VDDREF pch l=0.04u w=0.8u
m14852 578 425 VDDREF VDDREF pch l=0.04u w=0.8u
m14853 580 428 VDDREF VDDREF pch l=0.04u w=0.8u
m14854 581 429 VDDREF VDDREF pch l=0.04u w=0.8u
m14855 583 431 VDDREF VDDREF pch l=0.04u w=0.8u
m14856 584 432 VDDREF VDDREF pch l=0.04u w=0.8u
m14857 585 433 VDDREF VDDREF pch l=0.04u w=0.8u
m14858 587 435 VDDREF VDDREF pch l=0.04u w=0.8u
m14859 588 436 VDDREF VDDREF pch l=0.04u w=0.8u
m14860 VDDREF 559 564 VDDREF pch l=0.04u w=0.8u
m14861 589 550 VDDREF VDDREF pch l=0.04u w=0.8u
m14862 133 551 VDDREF VDDREF pch l=0.04u w=0.8u
m14863 590 552 VDDREF VDDREF pch l=0.04u w=0.8u
m14864 136 553 VDDREF VDDREF pch l=0.04u w=0.8u
m14865 591 554 VDDREF VDDREF pch l=0.04u w=0.8u
m14866 VDDREF 605 567 VDDREF pch l=0.04u w=0.8u
m14867 594 76 27633 VDDREF pch l=0.04u w=0.24u
m14868 592 555 VDDREF VDDREF pch l=0.04u w=0.8u
m14869 438 556 VDDREF VDDREF pch l=0.04u w=0.8u
m14870 VDDREF 606 VDDREF VDDREF pch l=0.26u w=1u
m14871 593 557 VDDREF VDDREF pch l=0.04u w=0.8u
m14872 442 558 VDDREF VDDREF pch l=0.04u w=0.8u
m14873 VDDREF 608 VDDREF VDDREF pch l=0.26u w=1u
m14874 568 206 393 VDDREF pch l=0.04u w=0.8u
m14875 477 610 571 VDDREF pch l=0.04u w=0.8u
m14876 569 209 394 VDDREF pch l=0.04u w=0.8u
m14877 597 611 574 VDDREF pch l=0.04u w=0.8u
m14878 599 612 577 VDDREF pch l=0.04u w=0.8u
m14879 600 613 579 VDDREF pch l=0.04u w=0.8u
m14880 62 614 582 VDDREF pch l=0.04u w=0.8u
m14881 64 615 586 VDDREF pch l=0.04u w=0.8u
m14882 VDDREF 617 VDDREF VDDREF pch l=0.26u w=1u
m14883 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14884 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14885 602 4328 548 VDDREF pch l=0.04u w=0.8u
m14886 603 4328 549 VDDREF pch l=0.04u w=0.8u
m14887 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m14888 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m14889 604 753 594 VDDREF pch l=0.04u w=0.8u
m14890 607 607 VDDREF VDDREF pch l=0.04u w=1u
m14891 609 609 VDDREF VDDREF pch l=0.04u w=1u
m14892 206 393 568 VDDREF pch l=0.04u w=0.8u
m14893 610 571 477 VDDREF pch l=0.04u w=0.8u
m14894 209 394 569 VDDREF pch l=0.04u w=0.8u
m14895 611 574 597 VDDREF pch l=0.04u w=0.8u
m14896 612 577 599 VDDREF pch l=0.04u w=0.8u
m14897 613 579 600 VDDREF pch l=0.04u w=0.8u
m14898 614 582 62 VDDREF pch l=0.04u w=0.8u
m14899 615 586 64 VDDREF pch l=0.04u w=0.8u
m14900 595 218 417 VDDREF pch l=0.04u w=0.8u
m14901 478 219 419 VDDREF pch l=0.04u w=0.8u
m14902 596 220 420 VDDREF pch l=0.04u w=0.8u
m14903 598 221 422 VDDREF pch l=0.04u w=0.8u
m14904 439 222 423 VDDREF pch l=0.04u w=0.8u
m14905 440 223 425 VDDREF pch l=0.04u w=0.8u
m14906 412 224 428 VDDREF pch l=0.04u w=0.8u
m14907 601 225 429 VDDREF pch l=0.04u w=0.8u
m14908 262 226 431 VDDREF pch l=0.04u w=0.8u
m14909 462 227 432 VDDREF pch l=0.04u w=0.8u
m14910 444 228 433 VDDREF pch l=0.04u w=0.8u
m14911 264 229 435 VDDREF pch l=0.04u w=0.8u
m14912 460 230 436 VDDREF pch l=0.04u w=0.8u
m14913 616 564 VDDREF VDDREF pch l=0.04u w=0.8u
m14914 618 618 VDDREF VDDREF pch l=0.04u w=1u
m14915 27653 565 602 VDDREF pch l=0.04u w=0.12u
m14916 27654 566 603 VDDREF pch l=0.04u w=0.12u
m14917 620 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14918 621 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14919 622 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14920 623 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m14921 619 520 591 VDDREF pch l=0.04u w=0.8u
m14922 605 652 VDDREF VDDREF pch l=0.04u w=0.8u
m14923 218 417 595 VDDREF pch l=0.04u w=0.8u
m14924 219 419 478 VDDREF pch l=0.04u w=0.8u
m14925 220 420 596 VDDREF pch l=0.04u w=0.8u
m14926 221 422 598 VDDREF pch l=0.04u w=0.8u
m14927 222 423 439 VDDREF pch l=0.04u w=0.8u
m14928 223 425 440 VDDREF pch l=0.04u w=0.8u
m14929 224 428 412 VDDREF pch l=0.04u w=0.8u
m14930 225 429 601 VDDREF pch l=0.04u w=0.8u
m14931 226 431 262 VDDREF pch l=0.04u w=0.8u
m14932 227 432 462 VDDREF pch l=0.04u w=0.8u
m14933 228 433 444 VDDREF pch l=0.04u w=0.8u
m14934 229 435 264 VDDREF pch l=0.04u w=0.8u
m14935 230 436 460 VDDREF pch l=0.04u w=0.8u
m14936 VDDREF 528 616 VDDREF pch l=0.04u w=0.8u
m14937 VDDREF 643 VDDREF VDDREF pch l=0.26u w=1u
m14938 VDDREF 644 VDDREF VDDREF pch l=0.26u w=1u
m14939 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m14940 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m14941 VDDREF 646 27653 VDDREF pch l=0.04u w=0.12u
m14942 VDDREF 647 27654 VDDREF pch l=0.04u w=0.12u
m14943 27668 76 619 VDDREF pch l=0.04u w=0.12u
m14944 VDDREF 2648 605 VDDREF pch l=0.04u w=0.8u
m14945 604 675 VDDREF VDDREF pch l=0.04u w=0.8u
m14946 635 710 VDDREF VDDREF pch l=0.04u w=0.8u
m14947 VDDREF 610 624 VDDREF pch l=0.04u w=0.8u
m14948 636 672 VDDREF VDDREF pch l=0.04u w=0.8u
m14949 VDDREF 611 625 VDDREF pch l=0.04u w=0.8u
m14950 VDDREF 612 626 VDDREF pch l=0.04u w=0.8u
m14951 VDDREF 613 627 VDDREF pch l=0.04u w=0.8u
m14952 VDDREF 614 628 VDDREF pch l=0.04u w=0.8u
m14953 VDDREF 615 629 VDDREF pch l=0.04u w=0.8u
m14954 VDDREF 630 631 VDDREF pch l=0.04u w=1u
m14955 642 642 VDDREF VDDREF pch l=0.04u w=1u
m14956 645 645 VDDREF VDDREF pch l=0.04u w=1u
m14957 646 602 VDDREF VDDREF pch l=0.04u w=0.8u
m14958 647 603 VDDREF VDDREF pch l=0.04u w=0.8u
m14959 VDDREF 259 27668 VDDREF pch l=0.04u w=0.12u
m14960 648 4328 633 VDDREF pch l=0.04u w=0.8u
m14961 649 4328 601 VDDREF pch l=0.04u w=0.8u
m14962 650 4328 634 VDDREF pch l=0.04u w=0.8u
m14963 651 4328 444 VDDREF pch l=0.04u w=0.8u
m14964 VDDREF 764 604 VDDREF pch l=0.04u w=0.8u
m14965 VDDREF 688 635 VDDREF pch l=0.04u w=0.8u
m14966 VDDREF 593 636 VDDREF pch l=0.04u w=0.8u
m14967 VDDREF 637 638 VDDREF pch l=0.04u w=1u
m14968 653 754 VDDREF VDDREF pch l=0.04u w=0.8u
m14969 654 736 VDDREF VDDREF pch l=0.04u w=0.8u
m14970 655 139 VDDREF VDDREF pch l=0.04u w=0.8u
m14971 656 755 VDDREF VDDREF pch l=0.04u w=0.8u
m14972 657 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m14973 658 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m14974 VDDREF 639 640 VDDREF pch l=0.04u w=1u
m14975 659 756 VDDREF VDDREF pch l=0.04u w=0.8u
m14976 660 FRAC[2] VDDREF VDDREF pch l=0.04u w=0.8u
m14977 VDDREF 704 641 VDDREF pch l=0.04u w=0.8u
m14978 661 737 VDDREF VDDREF pch l=0.04u w=0.8u
m14979 662 758 VDDREF VDDREF pch l=0.04u w=0.8u
m14980 663 634 VDDREF VDDREF pch l=0.04u w=0.8u
m14981 664 641 VDDREF VDDREF pch l=0.04u w=0.8u
m14982 665 756 VDDREF VDDREF pch l=0.04u w=0.8u
m14983 666 FRAC[2] VDDREF VDDREF pch l=0.04u w=0.8u
m14984 667 641 VDDREF VDDREF pch l=0.04u w=0.8u
m14985 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m14986 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m14987 259 619 VDDREF VDDREF pch l=0.04u w=0.8u
m14988 27714 620 648 VDDREF pch l=0.04u w=0.12u
m14989 27715 621 649 VDDREF pch l=0.04u w=0.12u
m14990 27716 622 650 VDDREF pch l=0.04u w=0.12u
m14991 27717 623 651 VDDREF pch l=0.04u w=0.12u
m14992 27719 604 VDDREF VDDREF pch l=0.04u w=0.12u
m14993 VDDREF 685 652 VDDREF pch l=0.04u w=0.8u
m14994 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m14995 VDDREF 731 653 VDDREF pch l=0.04u w=0.8u
m14996 274 823 VDDREF VDDREF pch l=0.04u w=0.8u
m14997 VDDREF 732 654 VDDREF pch l=0.04u w=0.8u
m14998 VDDREF 733 655 VDDREF pch l=0.04u w=0.8u
m14999 277 826 VDDREF VDDREF pch l=0.04u w=0.8u
m15000 VDDREF 734 656 VDDREF pch l=0.04u w=0.8u
m15001 VDDREF 893 657 VDDREF pch l=0.04u w=0.8u
m15002 VDDREF 894 658 VDDREF pch l=0.04u w=0.8u
m15003 VDDREF 735 659 VDDREF pch l=0.04u w=0.8u
m15004 280 829 VDDREF VDDREF pch l=0.04u w=0.8u
m15005 VDDREF 736 660 VDDREF pch l=0.04u w=0.8u
m15006 282 831 VDDREF VDDREF pch l=0.04u w=0.8u
m15007 VDDREF 131 661 VDDREF pch l=0.04u w=0.8u
m15008 VDDREF 737 662 VDDREF pch l=0.04u w=0.8u
m15009 285 834 VDDREF VDDREF pch l=0.04u w=0.8u
m15010 VDDREF 738 663 VDDREF pch l=0.04u w=0.8u
m15011 VDDREF 739 664 VDDREF pch l=0.04u w=0.8u
m15012 VDDREF 740 665 VDDREF pch l=0.04u w=0.8u
m15013 289 838 VDDREF VDDREF pch l=0.04u w=0.8u
m15014 VDDREF 741 666 VDDREF pch l=0.04u w=0.8u
m15015 VDDREF FBDIV[2] 667 VDDREF pch l=0.04u w=0.8u
m15016 VDDREF 669 668 VDDREF pch l=0.04u w=1u
m15017 VDDREF 670 671 VDDREF pch l=0.04u w=1u
m15018 673 565 646 VDDREF pch l=0.04u w=0.8u
m15019 674 566 647 VDDREF pch l=0.04u w=0.8u
m15020 VDDREF 679 27714 VDDREF pch l=0.04u w=0.12u
m15021 VDDREF 680 27715 VDDREF pch l=0.04u w=0.12u
m15022 VDDREF 681 27716 VDDREF pch l=0.04u w=0.12u
m15023 VDDREF 682 27717 VDDREF pch l=0.04u w=0.12u
m15024 675 753 27719 VDDREF pch l=0.04u w=0.12u
m15025 27876 567 VDDREF VDDREF pch l=0.04u w=0.24u
m15026 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15027 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15028 676 688 VDDREF VDDREF pch l=0.04u w=0.8u
m15029 VDDREF 712 274 VDDREF pch l=0.04u w=0.8u
m15030 677 593 VDDREF VDDREF pch l=0.04u w=0.8u
m15031 VDDREF 715 277 VDDREF pch l=0.04u w=0.8u
m15032 VDDREF 718 280 VDDREF pch l=0.04u w=0.8u
m15033 VDDREF 721 282 VDDREF pch l=0.04u w=0.8u
m15034 VDDREF 724 285 VDDREF pch l=0.04u w=0.8u
m15035 VDDREF 728 289 VDDREF pch l=0.04u w=0.8u
m15036 678 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15037 VDDREF 2197 672 VDDREF pch l=0.04u w=0.8u
m15038 VDDREF 705 VDDREF VDDREF pch l=0.26u w=1u
m15039 VDDREF 708 VDDREF VDDREF pch l=0.26u w=1u
m15040 28035 4328 673 VDDREF pch l=0.04u w=0.12u
m15041 28036 4328 674 VDDREF pch l=0.04u w=0.12u
m15042 679 648 VDDREF VDDREF pch l=0.04u w=0.8u
m15043 680 649 VDDREF VDDREF pch l=0.04u w=0.8u
m15044 681 650 VDDREF VDDREF pch l=0.04u w=0.8u
m15045 682 651 VDDREF VDDREF pch l=0.04u w=0.8u
m15046 683 259 VDDREF VDDREF pch l=0.04u w=0.8u
m15047 684 76 675 VDDREF pch l=0.04u w=0.8u
m15048 685 886 27876 VDDREF pch l=0.04u w=0.24u
m15049 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m15050 689 731 VDDREF VDDREF pch l=0.04u w=0.8u
m15051 690 732 VDDREF VDDREF pch l=0.04u w=0.8u
m15052 691 733 VDDREF VDDREF pch l=0.04u w=0.8u
m15053 692 734 VDDREF VDDREF pch l=0.04u w=0.8u
m15054 693 657 VDDREF VDDREF pch l=0.04u w=0.8u
m15055 694 658 VDDREF VDDREF pch l=0.04u w=0.8u
m15056 695 735 VDDREF VDDREF pch l=0.04u w=0.8u
m15057 696 736 VDDREF VDDREF pch l=0.04u w=0.8u
m15058 697 131 VDDREF VDDREF pch l=0.04u w=0.8u
m15059 698 737 VDDREF VDDREF pch l=0.04u w=0.8u
m15060 699 738 VDDREF VDDREF pch l=0.04u w=0.8u
m15061 700 739 VDDREF VDDREF pch l=0.04u w=0.8u
m15062 701 740 VDDREF VDDREF pch l=0.04u w=0.8u
m15063 702 741 VDDREF VDDREF pch l=0.04u w=0.8u
m15064 703 FBDIV[2] VDDREF VDDREF pch l=0.04u w=0.8u
m15065 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15066 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15067 706 706 VDDREF VDDREF pch l=0.04u w=1u
m15068 707 707 VDDREF VDDREF pch l=0.04u w=1u
m15069 VDDREF 747 28035 VDDREF pch l=0.04u w=0.12u
m15070 VDDREF 748 28036 VDDREF pch l=0.04u w=0.12u
m15071 VDDREF 259 683 VDDREF pch l=0.04u w=0.8u
m15072 709 847 685 VDDREF pch l=0.04u w=0.8u
m15073 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15074 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15075 686 710 688 VDDREF pch l=0.04u w=0.8u
m15076 712 571 VDDREF VDDREF pch l=0.04u w=0.8u
m15077 687 672 593 VDDREF pch l=0.04u w=0.8u
m15078 715 574 VDDREF VDDREF pch l=0.04u w=0.8u
m15079 718 577 VDDREF VDDREF pch l=0.04u w=0.8u
m15080 721 579 VDDREF VDDREF pch l=0.04u w=0.8u
m15081 724 582 VDDREF VDDREF pch l=0.04u w=0.8u
m15082 728 586 VDDREF VDDREF pch l=0.04u w=0.8u
m15083 720 4328 704 VDDREF pch l=0.04u w=0.8u
m15084 747 673 VDDREF VDDREF pch l=0.04u w=0.8u
m15085 748 674 VDDREF VDDREF pch l=0.04u w=0.8u
m15086 749 620 679 VDDREF pch l=0.04u w=0.8u
m15087 750 621 680 VDDREF pch l=0.04u w=0.8u
m15088 751 622 681 VDDREF pch l=0.04u w=0.8u
m15089 752 623 682 VDDREF pch l=0.04u w=0.8u
m15090 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m15091 753 76 VDDREF VDDREF pch l=0.04u w=0.8u
m15092 710 688 686 VDDREF pch l=0.04u w=0.8u
m15093 VDDREF 610 712 VDDREF pch l=0.04u w=0.8u
m15094 672 593 687 VDDREF pch l=0.04u w=0.8u
m15095 VDDREF 611 715 VDDREF pch l=0.04u w=0.8u
m15096 VDDREF 612 718 VDDREF pch l=0.04u w=0.8u
m15097 VDDREF 613 721 VDDREF pch l=0.04u w=0.8u
m15098 VDDREF 614 724 VDDREF pch l=0.04u w=0.8u
m15099 VDDREF 615 728 VDDREF pch l=0.04u w=0.8u
m15100 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15101 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15102 759 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15103 760 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15104 711 754 731 VDDREF pch l=0.04u w=0.8u
m15105 713 736 732 VDDREF pch l=0.04u w=0.8u
m15106 714 139 733 VDDREF pch l=0.04u w=0.8u
m15107 716 755 734 VDDREF pch l=0.04u w=0.8u
m15108 761 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15109 762 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15110 717 756 735 VDDREF pch l=0.04u w=0.8u
m15111 719 FRAC[2] 736 VDDREF pch l=0.04u w=0.8u
m15112 28057 678 720 VDDREF pch l=0.04u w=0.12u
m15113 722 737 131 VDDREF pch l=0.04u w=0.8u
m15114 723 758 737 VDDREF pch l=0.04u w=0.8u
m15115 725 634 738 VDDREF pch l=0.04u w=0.8u
m15116 726 641 739 VDDREF pch l=0.04u w=0.8u
m15117 727 756 740 VDDREF pch l=0.04u w=0.8u
m15118 729 FRAC[2] 741 VDDREF pch l=0.04u w=0.8u
m15119 730 641 FBDIV[2] VDDREF pch l=0.04u w=0.8u
m15120 VDDREF 743 744 VDDREF pch l=0.04u w=1u
m15121 VDDREF 746 745 VDDREF pch l=0.04u w=1u
m15122 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15123 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15124 28090 4328 749 VDDREF pch l=0.04u w=0.12u
m15125 28091 4328 750 VDDREF pch l=0.04u w=0.12u
m15126 28092 4328 751 VDDREF pch l=0.04u w=0.12u
m15127 28093 4328 752 VDDREF pch l=0.04u w=0.12u
m15128 763 683 VDDREF VDDREF pch l=0.04u w=0.8u
m15129 709 798 VDDREF VDDREF pch l=0.04u w=0.8u
m15130 754 731 711 VDDREF pch l=0.04u w=0.8u
m15131 736 732 713 VDDREF pch l=0.04u w=0.8u
m15132 139 733 714 VDDREF pch l=0.04u w=0.8u
m15133 755 734 716 VDDREF pch l=0.04u w=0.8u
m15134 756 735 717 VDDREF pch l=0.04u w=0.8u
m15135 FRAC[2] 736 719 VDDREF pch l=0.04u w=0.8u
m15136 VDDREF 778 28057 VDDREF pch l=0.04u w=0.12u
m15137 737 131 722 VDDREF pch l=0.04u w=0.8u
m15138 758 737 723 VDDREF pch l=0.04u w=0.8u
m15139 634 738 725 VDDREF pch l=0.04u w=0.8u
m15140 641 739 726 VDDREF pch l=0.04u w=0.8u
m15141 756 740 727 VDDREF pch l=0.04u w=0.8u
m15142 FRAC[2] 741 729 VDDREF pch l=0.04u w=0.8u
m15143 641 FBDIV[2] 730 VDDREF pch l=0.04u w=0.8u
m15144 771 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15145 772 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15146 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m15147 VDDREF 738 28090 VDDREF pch l=0.04u w=0.12u
m15148 VDDREF 443 28091 VDDREF pch l=0.04u w=0.12u
m15149 VDDREF 741 28092 VDDREF pch l=0.04u w=0.12u
m15150 VDDREF 445 28093 VDDREF pch l=0.04u w=0.12u
m15151 VDDREF 2648 709 VDDREF pch l=0.04u w=0.8u
m15152 VDDREF 236 764 VDDREF pch l=0.04u w=0.8u
m15153 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15154 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15155 765 686 VDDREF VDDREF pch l=0.04u w=0.8u
m15156 610 592 766 VDDREF pch l=0.04u w=0.8u
m15157 767 687 VDDREF VDDREF pch l=0.04u w=0.8u
m15158 611 599 139 VDDREF pch l=0.04u w=0.8u
m15159 612 593 FRAC[22] VDDREF pch l=0.04u w=0.8u
m15160 778 720 VDDREF VDDREF pch l=0.04u w=0.8u
m15161 613 793 202 VDDREF pch l=0.04u w=0.8u
m15162 614 202 64 VDDREF pch l=0.04u w=0.8u
m15163 615 204 FRAC[22] VDDREF pch l=0.04u w=0.8u
m15164 774 4328 769 VDDREF pch l=0.04u w=0.8u
m15165 775 4328 770 VDDREF pch l=0.04u w=0.8u
m15166 776 4328 693 VDDREF pch l=0.04u w=0.8u
m15167 777 4328 694 VDDREF pch l=0.04u w=0.8u
m15168 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15169 VDDREF 898 VDDREF VDDREF pch l=0.26u w=1u
m15170 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15171 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15172 738 749 VDDREF VDDREF pch l=0.04u w=0.8u
m15173 443 750 VDDREF VDDREF pch l=0.04u w=0.8u
m15174 741 751 VDDREF VDDREF pch l=0.04u w=0.8u
m15175 445 752 VDDREF VDDREF pch l=0.04u w=0.8u
m15176 792 763 VDDREF VDDREF pch l=0.04u w=0.8u
m15177 28410 709 VDDREF VDDREF pch l=0.04u w=0.12u
m15178 VDDREF 522 765 VDDREF pch l=0.04u w=0.8u
m15179 592 766 610 VDDREF pch l=0.04u w=0.8u
m15180 VDDREF 525 767 VDDREF pch l=0.04u w=0.8u
m15181 599 139 611 VDDREF pch l=0.04u w=0.8u
m15182 593 FRAC[22] 612 VDDREF pch l=0.04u w=0.8u
m15183 793 202 613 VDDREF pch l=0.04u w=0.8u
m15184 202 64 614 VDDREF pch l=0.04u w=0.8u
m15185 204 FRAC[22] 615 VDDREF pch l=0.04u w=0.8u
m15186 28415 759 774 VDDREF pch l=0.04u w=0.12u
m15187 28416 760 775 VDDREF pch l=0.04u w=0.12u
m15188 779 711 VDDREF VDDREF pch l=0.04u w=0.8u
m15189 780 713 VDDREF VDDREF pch l=0.04u w=0.8u
m15190 781 714 VDDREF VDDREF pch l=0.04u w=0.8u
m15191 782 716 VDDREF VDDREF pch l=0.04u w=0.8u
m15192 28417 761 776 VDDREF pch l=0.04u w=0.12u
m15193 28418 762 777 VDDREF pch l=0.04u w=0.12u
m15194 783 717 VDDREF VDDREF pch l=0.04u w=0.8u
m15195 784 719 VDDREF VDDREF pch l=0.04u w=0.8u
m15196 785 722 VDDREF VDDREF pch l=0.04u w=0.8u
m15197 786 723 VDDREF VDDREF pch l=0.04u w=0.8u
m15198 787 725 VDDREF VDDREF pch l=0.04u w=0.8u
m15199 788 726 VDDREF VDDREF pch l=0.04u w=0.8u
m15200 789 727 VDDREF VDDREF pch l=0.04u w=0.8u
m15201 790 729 VDDREF VDDREF pch l=0.04u w=0.8u
m15202 791 730 VDDREF VDDREF pch l=0.04u w=0.8u
m15203 794 155 VDDREF VDDREF pch l=0.04u w=0.8u
m15204 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m15205 795 4328 747 VDDREF pch l=0.04u w=0.8u
m15206 796 4328 748 VDDREF pch l=0.04u w=0.8u
m15207 797 810 792 VDDREF pch l=0.04u w=0.8u
m15208 798 847 28410 VDDREF pch l=0.04u w=0.12u
m15209 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15210 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15211 684 683 VDDREF VDDREF pch l=0.04u w=0.8u
m15212 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15213 VDDREF 898 VDDREF VDDREF pch l=0.26u w=1u
m15214 VDDREF 812 28415 VDDREF pch l=0.04u w=0.12u
m15215 VDDREF 813 28416 VDDREF pch l=0.04u w=0.12u
m15216 VDDREF 529 779 VDDREF pch l=0.04u w=0.8u
m15217 VDDREF 531 780 VDDREF pch l=0.04u w=0.8u
m15218 VDDREF 532 781 VDDREF pch l=0.04u w=0.8u
m15219 VDDREF 534 782 VDDREF pch l=0.04u w=0.8u
m15220 VDDREF 815 28417 VDDREF pch l=0.04u w=0.12u
m15221 VDDREF 816 28418 VDDREF pch l=0.04u w=0.12u
m15222 VDDREF 535 783 VDDREF pch l=0.04u w=0.8u
m15223 VDDREF 537 784 VDDREF pch l=0.04u w=0.8u
m15224 799 678 778 VDDREF pch l=0.04u w=0.8u
m15225 VDDREF 539 785 VDDREF pch l=0.04u w=0.8u
m15226 VDDREF 540 786 VDDREF pch l=0.04u w=0.8u
m15227 VDDREF 542 787 VDDREF pch l=0.04u w=0.8u
m15228 VDDREF 543 788 VDDREF pch l=0.04u w=0.8u
m15229 VDDREF 544 789 VDDREF pch l=0.04u w=0.8u
m15230 VDDREF 546 790 VDDREF pch l=0.04u w=0.8u
m15231 VDDREF 547 791 VDDREF pch l=0.04u w=0.8u
m15232 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15233 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15234 28483 771 795 VDDREF pch l=0.04u w=0.12u
m15235 28484 772 796 VDDREF pch l=0.04u w=0.12u
m15236 806 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15237 807 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15238 808 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15239 809 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15240 810 792 797 VDDREF pch l=0.04u w=0.8u
m15241 605 886 798 VDDREF pch l=0.04u w=0.8u
m15242 VDDREF 821 684 VDDREF pch l=0.04u w=0.8u
m15243 811 765 VDDREF VDDREF pch l=0.04u w=0.8u
m15244 812 774 VDDREF VDDREF pch l=0.04u w=0.8u
m15245 813 775 VDDREF VDDREF pch l=0.04u w=0.8u
m15246 VDDREF 592 800 VDDREF pch l=0.04u w=0.8u
m15247 814 767 VDDREF VDDREF pch l=0.04u w=0.8u
m15248 VDDREF 599 801 VDDREF pch l=0.04u w=0.8u
m15249 815 776 VDDREF VDDREF pch l=0.04u w=0.8u
m15250 816 777 VDDREF VDDREF pch l=0.04u w=0.8u
m15251 VDDREF 593 802 VDDREF pch l=0.04u w=0.8u
m15252 28491 4328 799 VDDREF pch l=0.04u w=0.12u
m15253 VDDREF 793 803 VDDREF pch l=0.04u w=0.8u
m15254 VDDREF 202 804 VDDREF pch l=0.04u w=0.8u
m15255 VDDREF 204 805 VDDREF pch l=0.04u w=0.8u
m15256 817 155 VDDREF VDDREF pch l=0.04u w=0.8u
m15257 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m15258 VDDREF 841 28483 VDDREF pch l=0.04u w=0.12u
m15259 VDDREF 842 28484 VDDREF pch l=0.04u w=0.12u
m15260 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15261 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15262 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15263 VDDREF 898 VDDREF VDDREF pch l=0.26u w=1u
m15264 VDDREF 635 811 VDDREF pch l=0.04u w=0.8u
m15265 VDDREF 636 814 VDDREF pch l=0.04u w=0.8u
m15266 VDDREF 852 28491 VDDREF pch l=0.04u w=0.12u
m15267 822 779 VDDREF VDDREF pch l=0.04u w=0.8u
m15268 824 780 VDDREF VDDREF pch l=0.04u w=0.8u
m15269 825 781 VDDREF VDDREF pch l=0.04u w=0.8u
m15270 827 782 VDDREF VDDREF pch l=0.04u w=0.8u
m15271 828 783 VDDREF VDDREF pch l=0.04u w=0.8u
m15272 830 784 VDDREF VDDREF pch l=0.04u w=0.8u
m15273 832 785 VDDREF VDDREF pch l=0.04u w=0.8u
m15274 833 786 VDDREF VDDREF pch l=0.04u w=0.8u
m15275 835 787 VDDREF VDDREF pch l=0.04u w=0.8u
m15276 836 788 VDDREF VDDREF pch l=0.04u w=0.8u
m15277 837 789 VDDREF VDDREF pch l=0.04u w=0.8u
m15278 839 790 VDDREF VDDREF pch l=0.04u w=0.8u
m15279 840 791 VDDREF VDDREF pch l=0.04u w=0.8u
m15280 VDDREF FBDIV[2] 817 VDDREF pch l=0.04u w=0.8u
m15281 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15282 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15283 841 795 VDDREF VDDREF pch l=0.04u w=0.8u
m15284 842 796 VDDREF VDDREF pch l=0.04u w=0.8u
m15285 843 4328 818 VDDREF pch l=0.04u w=0.8u
m15286 844 4328 819 VDDREF pch l=0.04u w=0.8u
m15287 845 4328 820 VDDREF pch l=0.04u w=0.8u
m15288 846 4328 739 VDDREF pch l=0.04u w=0.8u
m15289 847 886 VDDREF VDDREF pch l=0.04u w=0.8u
m15290 VDDREF 855 821 VDDREF pch l=0.04u w=0.8u
m15291 852 799 VDDREF VDDREF pch l=0.04u w=0.8u
m15292 848 759 812 VDDREF pch l=0.04u w=0.8u
m15293 849 760 813 VDDREF pch l=0.04u w=0.8u
m15294 VDDREF 653 822 VDDREF pch l=0.04u w=0.8u
m15295 823 592 VDDREF VDDREF pch l=0.04u w=0.8u
m15296 VDDREF 654 824 VDDREF pch l=0.04u w=0.8u
m15297 VDDREF 655 825 VDDREF pch l=0.04u w=0.8u
m15298 826 599 VDDREF VDDREF pch l=0.04u w=0.8u
m15299 VDDREF 656 827 VDDREF pch l=0.04u w=0.8u
m15300 850 761 815 VDDREF pch l=0.04u w=0.8u
m15301 851 762 816 VDDREF pch l=0.04u w=0.8u
m15302 VDDREF 659 828 VDDREF pch l=0.04u w=0.8u
m15303 829 593 VDDREF VDDREF pch l=0.04u w=0.8u
m15304 VDDREF 660 830 VDDREF pch l=0.04u w=0.8u
m15305 831 793 VDDREF VDDREF pch l=0.04u w=0.8u
m15306 VDDREF 661 832 VDDREF pch l=0.04u w=0.8u
m15307 VDDREF 662 833 VDDREF pch l=0.04u w=0.8u
m15308 834 202 VDDREF VDDREF pch l=0.04u w=0.8u
m15309 VDDREF 663 835 VDDREF pch l=0.04u w=0.8u
m15310 VDDREF 664 836 VDDREF pch l=0.04u w=0.8u
m15311 VDDREF 665 837 VDDREF pch l=0.04u w=0.8u
m15312 838 204 VDDREF VDDREF pch l=0.04u w=0.8u
m15313 VDDREF 666 839 VDDREF pch l=0.04u w=0.8u
m15314 VDDREF 667 840 VDDREF pch l=0.04u w=0.8u
m15315 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m15316 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15317 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15318 28507 806 843 VDDREF pch l=0.04u w=0.12u
m15319 28508 807 844 VDDREF pch l=0.04u w=0.12u
m15320 28509 808 845 VDDREF pch l=0.04u w=0.12u
m15321 28510 809 846 VDDREF pch l=0.04u w=0.12u
m15322 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15323 VDDREF 898 VDDREF VDDREF pch l=0.26u w=1u
m15324 853 377 VDDREF VDDREF pch l=0.04u w=0.8u
m15325 856 686 VDDREF VDDREF pch l=0.04u w=0.8u
m15326 28513 4328 848 VDDREF pch l=0.04u w=0.12u
m15327 28514 4328 849 VDDREF pch l=0.04u w=0.12u
m15328 VDDREF 766 823 VDDREF pch l=0.04u w=0.8u
m15329 857 687 VDDREF VDDREF pch l=0.04u w=0.8u
m15330 VDDREF 139 826 VDDREF pch l=0.04u w=0.8u
m15331 28515 4328 850 VDDREF pch l=0.04u w=0.12u
m15332 28516 4328 851 VDDREF pch l=0.04u w=0.12u
m15333 VDDREF FRAC[22] 829 VDDREF pch l=0.04u w=0.8u
m15334 VDDREF 202 831 VDDREF pch l=0.04u w=0.8u
m15335 VDDREF 64 834 VDDREF pch l=0.04u w=0.8u
m15336 VDDREF FRAC[22] 838 VDDREF pch l=0.04u w=0.8u
m15337 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15338 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15339 858 794 VDDREF VDDREF pch l=0.04u w=0.8u
m15340 859 771 841 VDDREF pch l=0.04u w=0.8u
m15341 860 772 842 VDDREF pch l=0.04u w=0.8u
m15342 VDDREF 881 28507 VDDREF pch l=0.04u w=0.12u
m15343 VDDREF 882 28508 VDDREF pch l=0.04u w=0.12u
m15344 VDDREF 883 28509 VDDREF pch l=0.04u w=0.12u
m15345 VDDREF 884 28510 VDDREF pch l=0.04u w=0.12u
m15346 VDDREF 886 854 VDDREF pch l=0.04u w=0.8u
m15347 VDDREF 1000 855 VDDREF pch l=0.04u w=0.8u
m15348 VDDREF 888 28513 VDDREF pch l=0.04u w=0.12u
m15349 VDDREF 732 28514 VDDREF pch l=0.04u w=0.12u
m15350 VDDREF 398 28515 VDDREF pch l=0.04u w=0.12u
m15351 VDDREF 736 28516 VDDREF pch l=0.04u w=0.12u
m15352 VDDREF 889 VDDREF VDDREF pch l=0.26u w=1u
m15353 862 711 VDDREF VDDREF pch l=0.04u w=0.8u
m15354 864 713 VDDREF VDDREF pch l=0.04u w=0.8u
m15355 865 714 VDDREF VDDREF pch l=0.04u w=0.8u
m15356 867 716 VDDREF VDDREF pch l=0.04u w=0.8u
m15357 868 717 VDDREF VDDREF pch l=0.04u w=0.8u
m15358 870 719 VDDREF VDDREF pch l=0.04u w=0.8u
m15359 872 722 VDDREF VDDREF pch l=0.04u w=0.8u
m15360 873 723 VDDREF VDDREF pch l=0.04u w=0.8u
m15361 875 725 VDDREF VDDREF pch l=0.04u w=0.8u
m15362 876 726 VDDREF VDDREF pch l=0.04u w=0.8u
m15363 877 727 VDDREF VDDREF pch l=0.04u w=0.8u
m15364 879 729 VDDREF VDDREF pch l=0.04u w=0.8u
m15365 880 730 VDDREF VDDREF pch l=0.04u w=0.8u
m15366 VDDREF 852 858 VDDREF pch l=0.04u w=0.8u
m15367 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15368 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15369 28526 4328 859 VDDREF pch l=0.04u w=0.12u
m15370 28527 4328 860 VDDREF pch l=0.04u w=0.12u
m15371 881 843 VDDREF VDDREF pch l=0.04u w=0.8u
m15372 882 844 VDDREF VDDREF pch l=0.04u w=0.8u
m15373 883 845 VDDREF VDDREF pch l=0.04u w=0.8u
m15374 884 846 VDDREF VDDREF pch l=0.04u w=0.8u
m15375 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15376 VDDREF 898 VDDREF VDDREF pch l=0.26u w=1u
m15377 885 377 VDDREF VDDREF pch l=0.04u w=0.8u
m15378 855 918 VDDREF VDDREF pch l=0.04u w=0.8u
m15379 888 848 VDDREF VDDREF pch l=0.04u w=0.8u
m15380 732 849 VDDREF VDDREF pch l=0.04u w=0.8u
m15381 VDDREF 899 VDDREF VDDREF pch l=0.26u w=1u
m15382 398 850 VDDREF VDDREF pch l=0.04u w=0.8u
m15383 736 851 VDDREF VDDREF pch l=0.04u w=0.8u
m15384 VDDREF 901 VDDREF VDDREF pch l=0.26u w=1u
m15385 890 890 VDDREF VDDREF pch l=0.04u w=1u
m15386 861 522 686 VDDREF pch l=0.04u w=0.8u
m15387 769 903 863 VDDREF pch l=0.04u w=0.8u
m15388 766 525 687 VDDREF pch l=0.04u w=0.8u
m15389 893 904 866 VDDREF pch l=0.04u w=0.8u
m15390 895 905 869 VDDREF pch l=0.04u w=0.8u
m15391 896 906 871 VDDREF pch l=0.04u w=0.8u
m15392 471 907 874 VDDREF pch l=0.04u w=0.8u
m15393 472 908 878 VDDREF pch l=0.04u w=0.8u
m15394 VDDREF 912 28526 VDDREF pch l=0.04u w=0.12u
m15395 VDDREF 913 28527 VDDREF pch l=0.04u w=0.12u
m15396 897 897 VDDREF VDDREF pch l=0.04u w=1u
m15397 VDDREF REFDIV[1] 885 VDDREF pch l=0.04u w=0.8u
m15398 886 930 VDDREF VDDREF pch l=0.04u w=0.8u
m15399 VDDREF 485 855 VDDREF pch l=0.04u w=0.8u
m15400 900 900 VDDREF VDDREF pch l=0.04u w=1u
m15401 902 902 VDDREF VDDREF pch l=0.04u w=1u
m15402 522 686 861 VDDREF pch l=0.04u w=0.8u
m15403 903 863 769 VDDREF pch l=0.04u w=0.8u
m15404 525 687 766 VDDREF pch l=0.04u w=0.8u
m15405 904 866 893 VDDREF pch l=0.04u w=0.8u
m15406 905 869 895 VDDREF pch l=0.04u w=0.8u
m15407 906 871 896 VDDREF pch l=0.04u w=0.8u
m15408 907 874 471 VDDREF pch l=0.04u w=0.8u
m15409 908 878 472 VDDREF pch l=0.04u w=0.8u
m15410 891 529 711 VDDREF pch l=0.04u w=0.8u
m15411 770 531 713 VDDREF pch l=0.04u w=0.8u
m15412 892 532 714 VDDREF pch l=0.04u w=0.8u
m15413 894 534 716 VDDREF pch l=0.04u w=0.8u
m15414 733 535 717 VDDREF pch l=0.04u w=0.8u
m15415 734 537 719 VDDREF pch l=0.04u w=0.8u
m15416 704 539 722 VDDREF pch l=0.04u w=0.8u
m15417 819 540 723 VDDREF pch l=0.04u w=0.8u
m15418 633 542 725 VDDREF pch l=0.04u w=0.8u
m15419 758 543 726 VDDREF pch l=0.04u w=0.8u
m15420 739 544 727 VDDREF pch l=0.04u w=0.8u
m15421 634 546 729 VDDREF pch l=0.04u w=0.8u
m15422 756 547 730 VDDREF pch l=0.04u w=0.8u
m15423 911 858 VDDREF VDDREF pch l=0.04u w=0.8u
m15424 VDDREF 926 VDDREF VDDREF pch l=0.26u w=1u
m15425 VDDREF 927 VDDREF VDDREF pch l=0.26u w=1u
m15426 912 859 VDDREF VDDREF pch l=0.04u w=0.8u
m15427 913 860 VDDREF VDDREF pch l=0.04u w=0.8u
m15428 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15429 914 806 881 VDDREF pch l=0.04u w=0.8u
m15430 915 807 882 VDDREF pch l=0.04u w=0.8u
m15431 916 808 883 VDDREF pch l=0.04u w=0.8u
m15432 917 809 884 VDDREF pch l=0.04u w=0.8u
m15433 VDDREF 2648 886 VDDREF pch l=0.04u w=0.8u
m15434 VDDREF 909 910 VDDREF pch l=0.04u w=1u
m15435 529 711 891 VDDREF pch l=0.04u w=0.8u
m15436 531 713 770 VDDREF pch l=0.04u w=0.8u
m15437 532 714 892 VDDREF pch l=0.04u w=0.8u
m15438 534 716 894 VDDREF pch l=0.04u w=0.8u
m15439 535 717 733 VDDREF pch l=0.04u w=0.8u
m15440 537 719 734 VDDREF pch l=0.04u w=0.8u
m15441 539 722 704 VDDREF pch l=0.04u w=0.8u
m15442 540 723 819 VDDREF pch l=0.04u w=0.8u
m15443 542 725 633 VDDREF pch l=0.04u w=0.8u
m15444 543 726 758 VDDREF pch l=0.04u w=0.8u
m15445 544 727 739 VDDREF pch l=0.04u w=0.8u
m15446 546 729 634 VDDREF pch l=0.04u w=0.8u
m15447 547 730 756 VDDREF pch l=0.04u w=0.8u
m15448 VDDREF 817 911 VDDREF pch l=0.04u w=0.8u
m15449 925 925 VDDREF VDDREF pch l=0.04u w=1u
m15450 928 928 VDDREF VDDREF pch l=0.04u w=1u
m15451 28556 4328 914 VDDREF pch l=0.04u w=0.12u
m15452 28557 4328 915 VDDREF pch l=0.04u w=0.12u
m15453 28558 4328 916 VDDREF pch l=0.04u w=0.12u
m15454 28559 4328 917 VDDREF pch l=0.04u w=0.12u
m15455 929 853 VDDREF VDDREF pch l=0.04u w=0.8u
m15456 VDDREF 944 918 VDDREF pch l=0.04u w=0.8u
m15457 931 1001 VDDREF VDDREF pch l=0.04u w=0.8u
m15458 VDDREF 903 919 VDDREF pch l=0.04u w=0.8u
m15459 932 962 VDDREF VDDREF pch l=0.04u w=0.8u
m15460 VDDREF 904 920 VDDREF pch l=0.04u w=0.8u
m15461 VDDREF 905 921 VDDREF pch l=0.04u w=0.8u
m15462 VDDREF 906 922 VDDREF pch l=0.04u w=0.8u
m15463 VDDREF 907 923 VDDREF pch l=0.04u w=0.8u
m15464 VDDREF 908 924 VDDREF pch l=0.04u w=0.8u
m15465 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15466 942 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15467 943 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15468 VDDREF 960 28556 VDDREF pch l=0.04u w=0.12u
m15469 VDDREF 737 28557 VDDREF pch l=0.04u w=0.12u
m15470 VDDREF 961 28558 VDDREF pch l=0.04u w=0.12u
m15471 VDDREF 740 28559 VDDREF pch l=0.04u w=0.12u
m15472 VDDREF 797 929 VDDREF pch l=0.04u w=0.8u
m15473 VDDREF 966 930 VDDREF pch l=0.04u w=0.8u
m15474 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15475 VDDREF 979 931 VDDREF pch l=0.04u w=0.8u
m15476 VDDREF 294 932 VDDREF pch l=0.04u w=0.8u
m15477 VDDREF 933 934 VDDREF pch l=0.04u w=1u
m15478 945 1041 VDDREF VDDREF pch l=0.04u w=0.8u
m15479 946 1028 VDDREF VDDREF pch l=0.04u w=0.8u
m15480 947 139 VDDREF VDDREF pch l=0.04u w=0.8u
m15481 948 1042 VDDREF VDDREF pch l=0.04u w=0.8u
m15482 949 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m15483 950 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m15484 VDDREF 935 936 VDDREF pch l=0.04u w=1u
m15485 951 1043 VDDREF VDDREF pch l=0.04u w=0.8u
m15486 952 FRAC[3] VDDREF VDDREF pch l=0.04u w=0.8u
m15487 VDDREF 995 937 VDDREF pch l=0.04u w=0.8u
m15488 953 1029 VDDREF VDDREF pch l=0.04u w=0.8u
m15489 954 1045 VDDREF VDDREF pch l=0.04u w=0.8u
m15490 955 998 VDDREF VDDREF pch l=0.04u w=0.8u
m15491 956 937 VDDREF VDDREF pch l=0.04u w=0.8u
m15492 957 1043 VDDREF VDDREF pch l=0.04u w=0.8u
m15493 958 FRAC[3] VDDREF VDDREF pch l=0.04u w=0.8u
m15494 959 937 VDDREF VDDREF pch l=0.04u w=0.8u
m15495 VDDREF 939 938 VDDREF pch l=0.04u w=1u
m15496 VDDREF 940 941 VDDREF pch l=0.04u w=1u
m15497 960 914 VDDREF VDDREF pch l=0.04u w=0.8u
m15498 737 915 VDDREF VDDREF pch l=0.04u w=0.8u
m15499 961 916 VDDREF VDDREF pch l=0.04u w=0.8u
m15500 740 917 VDDREF VDDREF pch l=0.04u w=0.8u
m15501 28579 854 VDDREF VDDREF pch l=0.04u w=0.24u
m15502 VDDREF 2194 944 VDDREF pch l=0.04u w=0.8u
m15503 VDDREF 1023 945 VDDREF pch l=0.04u w=0.8u
m15504 571 1114 VDDREF VDDREF pch l=0.04u w=0.8u
m15505 VDDREF 1024 946 VDDREF pch l=0.04u w=0.8u
m15506 VDDREF 1025 947 VDDREF pch l=0.04u w=0.8u
m15507 574 1117 VDDREF VDDREF pch l=0.04u w=0.8u
m15508 VDDREF 1026 948 VDDREF pch l=0.04u w=0.8u
m15509 VDDREF 1182 949 VDDREF pch l=0.04u w=0.8u
m15510 VDDREF 1183 950 VDDREF pch l=0.04u w=0.8u
m15511 VDDREF 1027 951 VDDREF pch l=0.04u w=0.8u
m15512 577 1120 VDDREF VDDREF pch l=0.04u w=0.8u
m15513 VDDREF 1028 952 VDDREF pch l=0.04u w=0.8u
m15514 579 1122 VDDREF VDDREF pch l=0.04u w=0.8u
m15515 VDDREF 131 953 VDDREF pch l=0.04u w=0.8u
m15516 VDDREF 1029 954 VDDREF pch l=0.04u w=0.8u
m15517 582 1125 VDDREF VDDREF pch l=0.04u w=0.8u
m15518 VDDREF 1030 955 VDDREF pch l=0.04u w=0.8u
m15519 VDDREF 999 956 VDDREF pch l=0.04u w=0.8u
m15520 VDDREF 1031 957 VDDREF pch l=0.04u w=0.8u
m15521 586 1129 VDDREF VDDREF pch l=0.04u w=0.8u
m15522 VDDREF 1032 958 VDDREF pch l=0.04u w=0.8u
m15523 VDDREF FBDIV[3] 959 VDDREF pch l=0.04u w=0.8u
m15524 VDDREF 970 VDDREF VDDREF pch l=0.26u w=1u
m15525 963 4328 912 VDDREF pch l=0.04u w=0.8u
m15526 964 4328 913 VDDREF pch l=0.04u w=0.8u
m15527 966 1152 28579 VDDREF pch l=0.04u w=0.24u
m15528 965 929 VDDREF VDDREF pch l=0.04u w=0.8u
m15529 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15530 944 1653 VDDREF VDDREF pch l=0.04u w=0.8u
m15531 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15532 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15533 967 979 VDDREF VDDREF pch l=0.04u w=0.8u
m15534 VDDREF 1004 571 VDDREF pch l=0.04u w=0.8u
m15535 968 294 VDDREF VDDREF pch l=0.04u w=0.8u
m15536 VDDREF 1007 574 VDDREF pch l=0.04u w=0.8u
m15537 VDDREF 1010 577 VDDREF pch l=0.04u w=0.8u
m15538 VDDREF 1013 579 VDDREF pch l=0.04u w=0.8u
m15539 VDDREF 1016 582 VDDREF pch l=0.04u w=0.8u
m15540 VDDREF 1020 586 VDDREF pch l=0.04u w=0.8u
m15541 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15542 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15543 969 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15544 971 971 VDDREF VDDREF pch l=0.04u w=1u
m15545 VDDREF 2465 962 VDDREF pch l=0.04u w=0.8u
m15546 28591 942 963 VDDREF pch l=0.04u w=0.12u
m15547 28592 943 964 VDDREF pch l=0.04u w=0.12u
m15548 972 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15549 973 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15550 974 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15551 975 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15552 976 1112 966 VDDREF pch l=0.04u w=0.8u
m15553 VDDREF 885 965 VDDREF pch l=0.04u w=0.8u
m15554 VDDREF 1061 944 VDDREF pch l=0.04u w=0.8u
m15555 980 1023 VDDREF VDDREF pch l=0.04u w=0.8u
m15556 981 1024 VDDREF VDDREF pch l=0.04u w=0.8u
m15557 982 1025 VDDREF VDDREF pch l=0.04u w=0.8u
m15558 983 1026 VDDREF VDDREF pch l=0.04u w=0.8u
m15559 984 949 VDDREF VDDREF pch l=0.04u w=0.8u
m15560 985 950 VDDREF VDDREF pch l=0.04u w=0.8u
m15561 986 1027 VDDREF VDDREF pch l=0.04u w=0.8u
m15562 987 1028 VDDREF VDDREF pch l=0.04u w=0.8u
m15563 988 131 VDDREF VDDREF pch l=0.04u w=0.8u
m15564 989 1029 VDDREF VDDREF pch l=0.04u w=0.8u
m15565 990 1030 VDDREF VDDREF pch l=0.04u w=0.8u
m15566 991 999 VDDREF VDDREF pch l=0.04u w=0.8u
m15567 992 1031 VDDREF VDDREF pch l=0.04u w=0.8u
m15568 993 1032 VDDREF VDDREF pch l=0.04u w=0.8u
m15569 994 FBDIV[3] VDDREF VDDREF pch l=0.04u w=0.8u
m15570 VDDREF 1035 28591 VDDREF pch l=0.04u w=0.12u
m15571 VDDREF 1036 28592 VDDREF pch l=0.04u w=0.12u
m15572 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15573 965 885 VDDREF VDDREF pch l=0.04u w=0.8u
m15574 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15575 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15576 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15577 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15578 977 1001 979 VDDREF pch l=0.04u w=0.8u
m15579 1004 863 VDDREF VDDREF pch l=0.04u w=0.8u
m15580 978 962 294 VDDREF pch l=0.04u w=0.8u
m15581 1007 866 VDDREF VDDREF pch l=0.04u w=0.8u
m15582 1010 869 VDDREF VDDREF pch l=0.04u w=0.8u
m15583 1013 871 VDDREF VDDREF pch l=0.04u w=0.8u
m15584 1016 874 VDDREF VDDREF pch l=0.04u w=0.8u
m15585 1020 878 VDDREF VDDREF pch l=0.04u w=0.8u
m15586 1012 4328 995 VDDREF pch l=0.04u w=0.8u
m15587 1035 963 VDDREF VDDREF pch l=0.04u w=0.8u
m15588 1036 964 VDDREF VDDREF pch l=0.04u w=0.8u
m15589 1037 4328 996 VDDREF pch l=0.04u w=0.8u
m15590 1038 4328 997 VDDREF pch l=0.04u w=0.8u
m15591 1039 4328 998 VDDREF pch l=0.04u w=0.8u
m15592 1040 4328 999 VDDREF pch l=0.04u w=0.8u
m15593 VDDREF 929 965 VDDREF pch l=0.04u w=0.8u
m15594 976 1085 VDDREF VDDREF pch l=0.04u w=0.8u
m15595 VDDREF 1240 1000 VDDREF pch l=0.04u w=0.8u
m15596 1001 979 977 VDDREF pch l=0.04u w=0.8u
m15597 VDDREF 903 1004 VDDREF pch l=0.04u w=0.8u
m15598 962 294 978 VDDREF pch l=0.04u w=0.8u
m15599 VDDREF 904 1007 VDDREF pch l=0.04u w=0.8u
m15600 VDDREF 905 1010 VDDREF pch l=0.04u w=0.8u
m15601 VDDREF 906 1013 VDDREF pch l=0.04u w=0.8u
m15602 VDDREF 907 1016 VDDREF pch l=0.04u w=0.8u
m15603 VDDREF 908 1020 VDDREF pch l=0.04u w=0.8u
m15604 1046 1055 VDDREF VDDREF pch l=0.04u w=0.8u
m15605 1047 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15606 1048 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15607 1003 1041 1023 VDDREF pch l=0.04u w=0.8u
m15608 1005 1028 1024 VDDREF pch l=0.04u w=0.8u
m15609 1006 139 1025 VDDREF pch l=0.04u w=0.8u
m15610 1008 1042 1026 VDDREF pch l=0.04u w=0.8u
m15611 1049 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15612 1050 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15613 1009 1043 1027 VDDREF pch l=0.04u w=0.8u
m15614 1011 FRAC[3] 1028 VDDREF pch l=0.04u w=0.8u
m15615 28614 969 1012 VDDREF pch l=0.04u w=0.12u
m15616 1014 1029 131 VDDREF pch l=0.04u w=0.8u
m15617 1015 1045 1029 VDDREF pch l=0.04u w=0.8u
m15618 1017 998 1030 VDDREF pch l=0.04u w=0.8u
m15619 1018 937 999 VDDREF pch l=0.04u w=0.8u
m15620 1019 1043 1031 VDDREF pch l=0.04u w=0.8u
m15621 1021 FRAC[3] 1032 VDDREF pch l=0.04u w=0.8u
m15622 1022 937 FBDIV[3] VDDREF pch l=0.04u w=0.8u
m15623 VDDREF 1080 1034 VDDREF pch l=0.04u w=0.8u
m15624 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15625 28618 972 1037 VDDREF pch l=0.04u w=0.12u
m15626 28619 973 1038 VDDREF pch l=0.04u w=0.12u
m15627 28620 974 1039 VDDREF pch l=0.04u w=0.12u
m15628 28621 975 1040 VDDREF pch l=0.04u w=0.12u
m15629 VDDREF 2648 976 VDDREF pch l=0.04u w=0.8u
m15630 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15631 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15632 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15633 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15634 1041 1023 1003 VDDREF pch l=0.04u w=0.8u
m15635 1028 1024 1005 VDDREF pch l=0.04u w=0.8u
m15636 139 1025 1006 VDDREF pch l=0.04u w=0.8u
m15637 1042 1026 1008 VDDREF pch l=0.04u w=0.8u
m15638 1043 1027 1009 VDDREF pch l=0.04u w=0.8u
m15639 FRAC[3] 1028 1011 VDDREF pch l=0.04u w=0.8u
m15640 VDDREF 1066 28614 VDDREF pch l=0.04u w=0.12u
m15641 1029 131 1014 VDDREF pch l=0.04u w=0.8u
m15642 1045 1029 1015 VDDREF pch l=0.04u w=0.8u
m15643 998 1030 1017 VDDREF pch l=0.04u w=0.8u
m15644 937 999 1018 VDDREF pch l=0.04u w=0.8u
m15645 1043 1031 1019 VDDREF pch l=0.04u w=0.8u
m15646 FRAC[3] 1032 1021 VDDREF pch l=0.04u w=0.8u
m15647 937 FBDIV[3] 1022 VDDREF pch l=0.04u w=0.8u
m15648 28623 1034 VDDREF VDDREF pch l=0.04u w=0.12u
m15649 1058 942 1035 VDDREF pch l=0.04u w=0.8u
m15650 1059 943 1036 VDDREF pch l=0.04u w=0.8u
m15651 VDDREF 1081 28618 VDDREF pch l=0.04u w=0.12u
m15652 VDDREF 1082 28619 VDDREF pch l=0.04u w=0.12u
m15653 VDDREF 1083 28620 VDDREF pch l=0.04u w=0.12u
m15654 VDDREF 1084 28621 VDDREF pch l=0.04u w=0.12u
m15655 28628 976 VDDREF VDDREF pch l=0.04u w=0.12u
m15656 1060 76 VDDREF VDDREF pch l=0.04u w=0.8u
m15657 1061 1090 VDDREF VDDREF pch l=0.04u w=0.8u
m15658 1052 977 VDDREF VDDREF pch l=0.04u w=0.8u
m15659 903 888 569 VDDREF pch l=0.04u w=0.8u
m15660 1053 978 VDDREF VDDREF pch l=0.04u w=0.8u
m15661 904 895 139 VDDREF pch l=0.04u w=0.8u
m15662 905 398 FRAC[21] VDDREF pch l=0.04u w=0.8u
m15663 1066 1012 VDDREF VDDREF pch l=0.04u w=0.8u
m15664 906 1086 589 VDDREF pch l=0.04u w=0.8u
m15665 907 589 472 VDDREF pch l=0.04u w=0.8u
m15666 908 590 FRAC[21] VDDREF pch l=0.04u w=0.8u
m15667 1051 1034 1055 VDDREF pch l=0.04u w=0.8u
m15668 1062 4328 1056 VDDREF pch l=0.04u w=0.8u
m15669 1063 4328 1057 VDDREF pch l=0.04u w=0.8u
m15670 1064 4328 984 VDDREF pch l=0.04u w=0.8u
m15671 1065 4328 985 VDDREF pch l=0.04u w=0.8u
m15672 1080 1593 28623 VDDREF pch l=0.04u w=0.12u
m15673 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15674 28636 4328 1058 VDDREF pch l=0.04u w=0.12u
m15675 28637 4328 1059 VDDREF pch l=0.04u w=0.12u
m15676 1081 1037 VDDREF VDDREF pch l=0.04u w=0.8u
m15677 1082 1038 VDDREF VDDREF pch l=0.04u w=0.8u
m15678 1083 1039 VDDREF VDDREF pch l=0.04u w=0.8u
m15679 1084 1040 VDDREF VDDREF pch l=0.04u w=0.8u
m15680 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15681 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15682 1085 1112 28628 VDDREF pch l=0.04u w=0.12u
m15683 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15684 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15685 VDDREF 1090 1061 VDDREF pch l=0.04u w=0.8u
m15686 VDDREF 811 1052 VDDREF pch l=0.04u w=0.8u
m15687 888 569 903 VDDREF pch l=0.04u w=0.8u
m15688 VDDREF 814 1053 VDDREF pch l=0.04u w=0.8u
m15689 895 139 904 VDDREF pch l=0.04u w=0.8u
m15690 398 FRAC[21] 905 VDDREF pch l=0.04u w=0.8u
m15691 1086 589 906 VDDREF pch l=0.04u w=0.8u
m15692 589 472 907 VDDREF pch l=0.04u w=0.8u
m15693 590 FRAC[21] 908 VDDREF pch l=0.04u w=0.8u
m15694 1034 1055 1051 VDDREF pch l=0.04u w=0.8u
m15695 28640 1047 1062 VDDREF pch l=0.04u w=0.12u
m15696 28641 1048 1063 VDDREF pch l=0.04u w=0.12u
m15697 1067 1003 VDDREF VDDREF pch l=0.04u w=0.8u
m15698 1068 1005 VDDREF VDDREF pch l=0.04u w=0.8u
m15699 1069 1006 VDDREF VDDREF pch l=0.04u w=0.8u
m15700 1070 1008 VDDREF VDDREF pch l=0.04u w=0.8u
m15701 28642 1049 1064 VDDREF pch l=0.04u w=0.12u
m15702 28643 1050 1065 VDDREF pch l=0.04u w=0.12u
m15703 1071 1009 VDDREF VDDREF pch l=0.04u w=0.8u
m15704 1072 1011 VDDREF VDDREF pch l=0.04u w=0.8u
m15705 1073 1014 VDDREF VDDREF pch l=0.04u w=0.8u
m15706 1074 1015 VDDREF VDDREF pch l=0.04u w=0.8u
m15707 1075 1017 VDDREF VDDREF pch l=0.04u w=0.8u
m15708 1076 1018 VDDREF VDDREF pch l=0.04u w=0.8u
m15709 1077 1019 VDDREF VDDREF pch l=0.04u w=0.8u
m15710 1078 1021 VDDREF VDDREF pch l=0.04u w=0.8u
m15711 1079 1022 VDDREF VDDREF pch l=0.04u w=0.8u
m15712 1087 1176 1080 VDDREF pch l=0.04u w=0.8u
m15713 1088 155 VDDREF VDDREF pch l=0.04u w=0.8u
m15714 VDDREF 1098 28636 VDDREF pch l=0.04u w=0.12u
m15715 VDDREF 1099 28637 VDDREF pch l=0.04u w=0.12u
m15716 886 1152 1085 VDDREF pch l=0.04u w=0.8u
m15717 1089 76 965 VDDREF pch l=0.04u w=0.8u
m15718 VDDREF 1105 28640 VDDREF pch l=0.04u w=0.12u
m15719 VDDREF 1106 28641 VDDREF pch l=0.04u w=0.12u
m15720 VDDREF 822 1067 VDDREF pch l=0.04u w=0.8u
m15721 VDDREF 824 1068 VDDREF pch l=0.04u w=0.8u
m15722 VDDREF 825 1069 VDDREF pch l=0.04u w=0.8u
m15723 VDDREF 827 1070 VDDREF pch l=0.04u w=0.8u
m15724 VDDREF 1108 28642 VDDREF pch l=0.04u w=0.12u
m15725 VDDREF 1109 28643 VDDREF pch l=0.04u w=0.12u
m15726 VDDREF 828 1071 VDDREF pch l=0.04u w=0.8u
m15727 VDDREF 830 1072 VDDREF pch l=0.04u w=0.8u
m15728 1091 969 1066 VDDREF pch l=0.04u w=0.8u
m15729 VDDREF 832 1073 VDDREF pch l=0.04u w=0.8u
m15730 VDDREF 833 1074 VDDREF pch l=0.04u w=0.8u
m15731 VDDREF 835 1075 VDDREF pch l=0.04u w=0.8u
m15732 VDDREF 836 1076 VDDREF pch l=0.04u w=0.8u
m15733 VDDREF 837 1077 VDDREF pch l=0.04u w=0.8u
m15734 VDDREF 839 1078 VDDREF pch l=0.04u w=0.8u
m15735 VDDREF 840 1079 VDDREF pch l=0.04u w=0.8u
m15736 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15737 1098 1058 VDDREF VDDREF pch l=0.04u w=0.8u
m15738 1099 1059 VDDREF VDDREF pch l=0.04u w=0.8u
m15739 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15740 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15741 1100 972 1081 VDDREF pch l=0.04u w=0.8u
m15742 1101 973 1082 VDDREF pch l=0.04u w=0.8u
m15743 1102 974 1083 VDDREF pch l=0.04u w=0.8u
m15744 1103 975 1084 VDDREF pch l=0.04u w=0.8u
m15745 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15746 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15747 28652 1060 1089 VDDREF pch l=0.04u w=0.12u
m15748 VDDREF 1137 1090 VDDREF pch l=0.04u w=0.8u
m15749 1104 1052 VDDREF VDDREF pch l=0.04u w=0.8u
m15750 1105 1062 VDDREF VDDREF pch l=0.04u w=0.8u
m15751 1106 1063 VDDREF VDDREF pch l=0.04u w=0.8u
m15752 VDDREF 888 1092 VDDREF pch l=0.04u w=0.8u
m15753 1107 1053 VDDREF VDDREF pch l=0.04u w=0.8u
m15754 VDDREF 895 1093 VDDREF pch l=0.04u w=0.8u
m15755 1108 1064 VDDREF VDDREF pch l=0.04u w=0.8u
m15756 1109 1065 VDDREF VDDREF pch l=0.04u w=0.8u
m15757 VDDREF 398 1094 VDDREF pch l=0.04u w=0.8u
m15758 28653 4328 1091 VDDREF pch l=0.04u w=0.12u
m15759 VDDREF 1086 1095 VDDREF pch l=0.04u w=0.8u
m15760 VDDREF 589 1096 VDDREF pch l=0.04u w=0.8u
m15761 VDDREF 590 1097 VDDREF pch l=0.04u w=0.8u
m15762 1110 PD VDDREF VDDREF pch l=0.04u w=0.8u
m15763 VDDREF 1143 1087 VDDREF pch l=0.04u w=0.8u
m15764 1111 155 VDDREF VDDREF pch l=0.04u w=0.8u
m15765 28658 4328 1100 VDDREF pch l=0.04u w=0.12u
m15766 28659 4328 1101 VDDREF pch l=0.04u w=0.12u
m15767 28660 4328 1102 VDDREF pch l=0.04u w=0.12u
m15768 28661 4328 1103 VDDREF pch l=0.04u w=0.12u
m15769 1112 1152 VDDREF VDDREF pch l=0.04u w=0.8u
m15770 VDDREF 1135 28652 VDDREF pch l=0.04u w=0.12u
m15771 28663 1090 VDDREF VDDREF pch l=0.04u w=0.12u
m15772 VDDREF 931 1104 VDDREF pch l=0.04u w=0.8u
m15773 VDDREF 932 1107 VDDREF pch l=0.04u w=0.8u
m15774 VDDREF 1142 28653 VDDREF pch l=0.04u w=0.12u
m15775 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15776 1113 1067 VDDREF VDDREF pch l=0.04u w=0.8u
m15777 1115 1068 VDDREF VDDREF pch l=0.04u w=0.8u
m15778 1116 1069 VDDREF VDDREF pch l=0.04u w=0.8u
m15779 1118 1070 VDDREF VDDREF pch l=0.04u w=0.8u
m15780 1119 1071 VDDREF VDDREF pch l=0.04u w=0.8u
m15781 1121 1072 VDDREF VDDREF pch l=0.04u w=0.8u
m15782 1123 1073 VDDREF VDDREF pch l=0.04u w=0.8u
m15783 1124 1074 VDDREF VDDREF pch l=0.04u w=0.8u
m15784 1126 1075 VDDREF VDDREF pch l=0.04u w=0.8u
m15785 1127 1076 VDDREF VDDREF pch l=0.04u w=0.8u
m15786 1128 1077 VDDREF VDDREF pch l=0.04u w=0.8u
m15787 1130 1078 VDDREF VDDREF pch l=0.04u w=0.8u
m15788 1131 1079 VDDREF VDDREF pch l=0.04u w=0.8u
m15789 28669 1087 VDDREF VDDREF pch l=0.04u w=0.12u
m15790 VDDREF FBDIV[3] 1111 VDDREF pch l=0.04u w=0.8u
m15791 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15792 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15793 1133 1146 VDDREF VDDREF pch l=0.04u w=0.8u
m15794 1134 70 VDDREF VDDREF pch l=0.04u w=0.8u
m15795 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15796 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15797 VDDREF 1030 28658 VDDREF pch l=0.04u w=0.12u
m15798 VDDREF 1029 28659 VDDREF pch l=0.04u w=0.12u
m15799 VDDREF 1032 28660 VDDREF pch l=0.04u w=0.12u
m15800 VDDREF 1031 28661 VDDREF pch l=0.04u w=0.12u
m15801 1135 1089 VDDREF VDDREF pch l=0.04u w=0.8u
m15802 1137 76 28663 VDDREF pch l=0.04u w=0.12u
m15803 1142 1091 VDDREF VDDREF pch l=0.04u w=0.8u
m15804 1138 1047 1105 VDDREF pch l=0.04u w=0.8u
m15805 1139 1048 1106 VDDREF pch l=0.04u w=0.8u
m15806 VDDREF 945 1113 VDDREF pch l=0.04u w=0.8u
m15807 1114 888 VDDREF VDDREF pch l=0.04u w=0.8u
m15808 VDDREF 946 1115 VDDREF pch l=0.04u w=0.8u
m15809 VDDREF 947 1116 VDDREF pch l=0.04u w=0.8u
m15810 1117 895 VDDREF VDDREF pch l=0.04u w=0.8u
m15811 VDDREF 948 1118 VDDREF pch l=0.04u w=0.8u
m15812 1140 1049 1108 VDDREF pch l=0.04u w=0.8u
m15813 1141 1050 1109 VDDREF pch l=0.04u w=0.8u
m15814 VDDREF 951 1119 VDDREF pch l=0.04u w=0.8u
m15815 1120 398 VDDREF VDDREF pch l=0.04u w=0.8u
m15816 VDDREF 952 1121 VDDREF pch l=0.04u w=0.8u
m15817 1122 1086 VDDREF VDDREF pch l=0.04u w=0.8u
m15818 VDDREF 953 1123 VDDREF pch l=0.04u w=0.8u
m15819 VDDREF 954 1124 VDDREF pch l=0.04u w=0.8u
m15820 1125 589 VDDREF VDDREF pch l=0.04u w=0.8u
m15821 VDDREF 955 1126 VDDREF pch l=0.04u w=0.8u
m15822 VDDREF 956 1127 VDDREF pch l=0.04u w=0.8u
m15823 VDDREF 957 1128 VDDREF pch l=0.04u w=0.8u
m15824 1129 590 VDDREF VDDREF pch l=0.04u w=0.8u
m15825 VDDREF 958 1130 VDDREF pch l=0.04u w=0.8u
m15826 VDDREF 959 1131 VDDREF pch l=0.04u w=0.8u
m15827 1143 1176 28669 VDDREF pch l=0.04u w=0.12u
m15828 VDDREF 1372 1132 VDDREF pch l=0.04u w=0.8u
m15829 1030 1100 VDDREF VDDREF pch l=0.04u w=0.8u
m15830 1029 1101 VDDREF VDDREF pch l=0.04u w=0.8u
m15831 1032 1102 VDDREF VDDREF pch l=0.04u w=0.8u
m15832 1031 1103 VDDREF VDDREF pch l=0.04u w=0.8u
m15833 VDDREF 1152 1136 VDDREF pch l=0.04u w=0.8u
m15834 1147 1241 1137 VDDREF pch l=0.04u w=0.8u
m15835 VDDREF 1153 VDDREF VDDREF pch l=0.26u w=1u
m15836 1148 977 VDDREF VDDREF pch l=0.04u w=0.8u
m15837 28680 4328 1138 VDDREF pch l=0.04u w=0.12u
m15838 28681 4328 1139 VDDREF pch l=0.04u w=0.12u
m15839 VDDREF 569 1114 VDDREF pch l=0.04u w=0.8u
m15840 1149 978 VDDREF VDDREF pch l=0.04u w=0.8u
m15841 VDDREF 139 1117 VDDREF pch l=0.04u w=0.8u
m15842 28682 4328 1140 VDDREF pch l=0.04u w=0.12u
m15843 28683 4328 1141 VDDREF pch l=0.04u w=0.12u
m15844 VDDREF FRAC[21] 1120 VDDREF pch l=0.04u w=0.8u
m15845 VDDREF 589 1122 VDDREF pch l=0.04u w=0.8u
m15846 VDDREF 472 1125 VDDREF pch l=0.04u w=0.8u
m15847 VDDREF FRAC[21] 1129 VDDREF pch l=0.04u w=0.8u
m15848 1055 1593 1143 VDDREF pch l=0.04u w=0.8u
m15849 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15850 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15851 1150 1088 VDDREF VDDREF pch l=0.04u w=0.8u
m15852 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15853 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15854 1144 1098 1146 VDDREF pch l=0.04u w=0.8u
m15855 1145 1099 70 VDDREF pch l=0.04u w=0.8u
m15856 1151 1060 1135 VDDREF pch l=0.04u w=0.8u
m15857 1154 1154 VDDREF VDDREF pch l=0.04u w=1u
m15858 VDDREF 1179 28680 VDDREF pch l=0.04u w=0.12u
m15859 VDDREF 1024 28681 VDDREF pch l=0.04u w=0.12u
m15860 VDDREF 94 28682 VDDREF pch l=0.04u w=0.12u
m15861 VDDREF 1028 28683 VDDREF pch l=0.04u w=0.12u
m15862 318 1156 VDDREF VDDREF pch l=0.04u w=0.8u
m15863 1158 1003 VDDREF VDDREF pch l=0.04u w=0.8u
m15864 1160 1005 VDDREF VDDREF pch l=0.04u w=0.8u
m15865 1161 1006 VDDREF VDDREF pch l=0.04u w=0.8u
m15866 1163 1008 VDDREF VDDREF pch l=0.04u w=0.8u
m15867 1164 1009 VDDREF VDDREF pch l=0.04u w=0.8u
m15868 1166 1011 VDDREF VDDREF pch l=0.04u w=0.8u
m15869 1167 1014 VDDREF VDDREF pch l=0.04u w=0.8u
m15870 1168 1015 VDDREF VDDREF pch l=0.04u w=0.8u
m15871 1170 1017 VDDREF VDDREF pch l=0.04u w=0.8u
m15872 1171 1018 VDDREF VDDREF pch l=0.04u w=0.8u
m15873 1172 1019 VDDREF VDDREF pch l=0.04u w=0.8u
m15874 1174 1021 VDDREF VDDREF pch l=0.04u w=0.8u
m15875 1175 1022 VDDREF VDDREF pch l=0.04u w=0.8u
m15876 1157 1372 1051 VDDREF pch l=0.04u w=0.8u
m15877 VDDREF 1142 1150 VDDREF pch l=0.04u w=0.8u
m15878 1098 1146 1144 VDDREF pch l=0.04u w=0.8u
m15879 1099 70 1145 VDDREF pch l=0.04u w=0.8u
m15880 28696 76 1151 VDDREF pch l=0.04u w=0.12u
m15881 1152 1201 VDDREF VDDREF pch l=0.04u w=0.8u
m15882 VDDREF 1202 1147 VDDREF pch l=0.04u w=0.8u
m15883 1179 1138 VDDREF VDDREF pch l=0.04u w=0.8u
m15884 1024 1139 VDDREF VDDREF pch l=0.04u w=0.8u
m15885 VDDREF 1186 VDDREF VDDREF pch l=0.26u w=1u
m15886 94 1140 VDDREF VDDREF pch l=0.04u w=0.8u
m15887 1028 1141 VDDREF VDDREF pch l=0.04u w=0.8u
m15888 VDDREF 1188 VDDREF VDDREF pch l=0.26u w=1u
m15889 1155 811 977 VDDREF pch l=0.04u w=0.8u
m15890 1056 1190 1159 VDDREF pch l=0.04u w=0.8u
m15891 474 814 978 VDDREF pch l=0.04u w=0.8u
m15892 1182 1191 1162 VDDREF pch l=0.04u w=0.8u
m15893 1184 1192 1165 VDDREF pch l=0.04u w=0.8u
m15894 1185 1193 131 VDDREF pch l=0.04u w=0.8u
m15895 818 1194 1169 VDDREF pch l=0.04u w=0.8u
m15896 820 1195 1173 VDDREF pch l=0.04u w=0.8u
m15897 VDDREF 1593 1176 VDDREF pch l=0.04u w=0.8u
m15898 28702 1132 1157 VDDREF pch l=0.04u w=0.12u
m15899 VDDREF 1197 VDDREF VDDREF pch l=0.26u w=1u
m15900 VDDREF 1198 VDDREF VDDREF pch l=0.26u w=1u
m15901 VDDREF 810 28696 VDDREF pch l=0.04u w=0.12u
m15902 VDDREF 2648 1152 VDDREF pch l=0.04u w=0.8u
m15903 28706 1147 VDDREF VDDREF pch l=0.04u w=0.12u
m15904 VDDREF 1177 1178 VDDREF pch l=0.04u w=1u
m15905 1187 1187 VDDREF VDDREF pch l=0.04u w=1u
m15906 1189 1189 VDDREF VDDREF pch l=0.04u w=1u
m15907 811 977 1155 VDDREF pch l=0.04u w=0.8u
m15908 1190 1159 1056 VDDREF pch l=0.04u w=0.8u
m15909 814 978 474 VDDREF pch l=0.04u w=0.8u
m15910 1191 1162 1182 VDDREF pch l=0.04u w=0.8u
m15911 1192 1165 1184 VDDREF pch l=0.04u w=0.8u
m15912 1193 131 1185 VDDREF pch l=0.04u w=0.8u
m15913 1194 1169 818 VDDREF pch l=0.04u w=0.8u
m15914 1195 1173 820 VDDREF pch l=0.04u w=0.8u
m15915 VDDREF 1204 28702 VDDREF pch l=0.04u w=0.12u
m15916 1196 1196 VDDREF VDDREF pch l=0.04u w=1u
m15917 1199 1199 VDDREF VDDREF pch l=0.04u w=1u
m15918 1180 822 1003 VDDREF pch l=0.04u w=0.8u
m15919 1057 824 1005 VDDREF pch l=0.04u w=0.8u
m15920 1181 825 1006 VDDREF pch l=0.04u w=0.8u
m15921 1183 827 1008 VDDREF pch l=0.04u w=0.8u
m15922 1025 828 1009 VDDREF pch l=0.04u w=0.8u
m15923 1026 830 1011 VDDREF pch l=0.04u w=0.8u
m15924 995 832 1014 VDDREF pch l=0.04u w=0.8u
m15925 997 833 1015 VDDREF pch l=0.04u w=0.8u
m15926 996 835 1017 VDDREF pch l=0.04u w=0.8u
m15927 1045 836 1018 VDDREF pch l=0.04u w=0.8u
m15928 999 837 1019 VDDREF pch l=0.04u w=0.8u
m15929 998 839 1021 VDDREF pch l=0.04u w=0.8u
m15930 1043 840 1022 VDDREF pch l=0.04u w=0.8u
m15931 1200 1150 VDDREF VDDREF pch l=0.04u w=0.8u
m15932 810 1151 VDDREF VDDREF pch l=0.04u w=0.8u
m15933 1202 1241 28706 VDDREF pch l=0.04u w=0.12u
m15934 1203 1203 VDDREF VDDREF pch l=0.04u w=1u
m15935 1204 1110 VDDREF VDDREF pch l=0.04u w=0.8u
m15936 822 1003 1180 VDDREF pch l=0.04u w=0.8u
m15937 824 1005 1057 VDDREF pch l=0.04u w=0.8u
m15938 825 1006 1181 VDDREF pch l=0.04u w=0.8u
m15939 827 1008 1183 VDDREF pch l=0.04u w=0.8u
m15940 828 1009 1025 VDDREF pch l=0.04u w=0.8u
m15941 830 1011 1026 VDDREF pch l=0.04u w=0.8u
m15942 832 1014 995 VDDREF pch l=0.04u w=0.8u
m15943 833 1015 997 VDDREF pch l=0.04u w=0.8u
m15944 835 1017 996 VDDREF pch l=0.04u w=0.8u
m15945 836 1018 1045 VDDREF pch l=0.04u w=0.8u
m15946 837 1019 999 VDDREF pch l=0.04u w=0.8u
m15947 839 1021 998 VDDREF pch l=0.04u w=0.8u
m15948 840 1022 1043 VDDREF pch l=0.04u w=0.8u
m15949 VDDREF 1257 1055 VDDREF pch l=0.04u w=0.8u
m15950 VDDREF 1111 1200 VDDREF pch l=0.04u w=0.8u
m15951 1223 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15952 1224 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m15953 VDDREF 1258 1201 VDDREF pch l=0.04u w=0.8u
m15954 1225 76 1202 VDDREF pch l=0.04u w=0.8u
m15955 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m15956 VDDREF 1157 1204 VDDREF pch l=0.04u w=0.8u
m15957 1226 1104 VDDREF VDDREF pch l=0.04u w=0.8u
m15958 VDDREF 1190 1205 VDDREF pch l=0.04u w=0.8u
m15959 1227 1107 VDDREF VDDREF pch l=0.04u w=0.8u
m15960 VDDREF 1191 1206 VDDREF pch l=0.04u w=0.8u
m15961 VDDREF 1192 1207 VDDREF pch l=0.04u w=0.8u
m15962 VDDREF 1193 1208 VDDREF pch l=0.04u w=0.8u
m15963 VDDREF 1210 1209 VDDREF pch l=0.04u w=1u
m15964 VDDREF 1211 1212 VDDREF pch l=0.04u w=1u
m15965 VDDREF 1194 1213 VDDREF pch l=0.04u w=0.8u
m15966 VDDREF 1215 1214 VDDREF pch l=0.04u w=1u
m15967 VDDREF 1216 1217 VDDREF pch l=0.04u w=1u
m15968 VDDREF 1195 1218 VDDREF pch l=0.04u w=0.8u
m15969 28730 1055 VDDREF VDDREF pch l=0.04u w=0.12u
m15970 VDDREF 1220 1219 VDDREF pch l=0.04u w=1u
m15971 VDDREF 1221 1222 VDDREF pch l=0.04u w=1u
m15972 1240 810 VDDREF VDDREF pch l=0.04u w=0.8u
m15973 28732 1136 VDDREF VDDREF pch l=0.04u w=0.24u
m15974 1257 1372 28730 VDDREF pch l=0.04u w=0.12u
m15975 1242 1113 VDDREF VDDREF pch l=0.04u w=0.8u
m15976 1243 1115 VDDREF VDDREF pch l=0.04u w=0.8u
m15977 1244 1116 VDDREF VDDREF pch l=0.04u w=0.8u
m15978 1245 1118 VDDREF VDDREF pch l=0.04u w=0.8u
m15979 1246 1119 VDDREF VDDREF pch l=0.04u w=0.8u
m15980 1247 1121 VDDREF VDDREF pch l=0.04u w=0.8u
m15981 1250 1123 VDDREF VDDREF pch l=0.04u w=0.8u
m15982 1251 1124 VDDREF VDDREF pch l=0.04u w=0.8u
m15983 1252 1126 VDDREF VDDREF pch l=0.04u w=0.8u
m15984 1253 1127 VDDREF VDDREF pch l=0.04u w=0.8u
m15985 1254 1128 VDDREF VDDREF pch l=0.04u w=0.8u
m15986 1255 1130 VDDREF VDDREF pch l=0.04u w=0.8u
m15987 1256 1131 VDDREF VDDREF pch l=0.04u w=0.8u
m15988 1248 4328 1144 VDDREF pch l=0.04u w=0.8u
m15989 1249 4328 1145 VDDREF pch l=0.04u w=0.8u
m15990 VDDREF 1228 1229 VDDREF pch l=0.04u w=1u
m15991 VDDREF 1231 1230 VDDREF pch l=0.04u w=1u
m15992 VDDREF 1232 1233 VDDREF pch l=0.04u w=1u
m15993 VDDREF 1234 1235 VDDREF pch l=0.04u w=1u
m15994 VDDREF 1237 1236 VDDREF pch l=0.04u w=1u
m15995 VDDREF 1238 1239 VDDREF pch l=0.04u w=1u
m15996 VDDREF 810 1240 VDDREF pch l=0.04u w=0.8u
m15997 1258 1392 28732 VDDREF pch l=0.04u w=0.24u
m15998 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m15999 VDDREF 76 1241 VDDREF pch l=0.04u w=0.8u
m16000 VDDREF 1346 VDDREF VDDREF pch l=0.26u w=1u
m16001 VDDREF 1347 VDDREF VDDREF pch l=0.26u w=1u
m16002 VDDREF 1350 VDDREF VDDREF pch l=0.26u w=1u
m16003 VDDREF 1351 VDDREF VDDREF pch l=0.26u w=1u
m16004 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16005 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16006 1260 1315 1257 VDDREF pch l=0.04u w=0.8u
m16007 1259 1132 1204 VDDREF pch l=0.04u w=0.8u
m16008 1261 89 VDDREF VDDREF pch l=0.04u w=0.8u
m16009 863 1373 VDDREF VDDREF pch l=0.04u w=0.8u
m16010 1262 90 VDDREF VDDREF pch l=0.04u w=0.8u
m16011 866 1374 VDDREF VDDREF pch l=0.04u w=0.8u
m16012 869 1375 VDDREF VDDREF pch l=0.04u w=0.8u
m16013 871 1376 VDDREF VDDREF pch l=0.04u w=0.8u
m16014 874 1377 VDDREF VDDREF pch l=0.04u w=0.8u
m16015 878 1378 VDDREF VDDREF pch l=0.04u w=0.8u
m16016 28749 1223 1248 VDDREF pch l=0.04u w=0.12u
m16017 28750 1224 1249 VDDREF pch l=0.04u w=0.12u
m16018 1266 1353 1258 VDDREF pch l=0.04u w=0.8u
m16019 28756 1372 1259 VDDREF pch l=0.04u w=0.24u
m16020 VDDREF 393 1261 VDDREF pch l=0.04u w=0.8u
m16021 VDDREF 1284 863 VDDREF pch l=0.04u w=0.8u
m16022 VDDREF 394 1262 VDDREF pch l=0.04u w=0.8u
m16023 VDDREF 1285 866 VDDREF pch l=0.04u w=0.8u
m16024 VDDREF 1286 869 VDDREF pch l=0.04u w=0.8u
m16025 VDDREF 1287 871 VDDREF pch l=0.04u w=0.8u
m16026 VDDREF 1288 874 VDDREF pch l=0.04u w=0.8u
m16027 VDDREF 1289 878 VDDREF pch l=0.04u w=0.8u
m16028 1267 111 VDDREF VDDREF pch l=0.04u w=0.8u
m16029 1268 112 VDDREF VDDREF pch l=0.04u w=0.8u
m16030 1269 113 VDDREF VDDREF pch l=0.04u w=0.8u
m16031 1270 114 VDDREF VDDREF pch l=0.04u w=0.8u
m16032 1271 115 VDDREF VDDREF pch l=0.04u w=0.8u
m16033 1272 116 VDDREF VDDREF pch l=0.04u w=0.8u
m16034 VDDREF 1281 28749 VDDREF pch l=0.04u w=0.12u
m16035 VDDREF 1282 28750 VDDREF pch l=0.04u w=0.12u
m16036 1273 118 VDDREF VDDREF pch l=0.04u w=0.8u
m16037 1274 119 VDDREF VDDREF pch l=0.04u w=0.8u
m16038 1275 120 VDDREF VDDREF pch l=0.04u w=0.8u
m16039 1276 121 VDDREF VDDREF pch l=0.04u w=0.8u
m16040 1277 122 VDDREF VDDREF pch l=0.04u w=0.8u
m16041 1278 123 VDDREF VDDREF pch l=0.04u w=0.8u
m16042 1279 124 VDDREF VDDREF pch l=0.04u w=0.8u
m16043 VDDREF 1265 1264 VDDREF pch l=0.04u w=1u
m16044 VDDREF 1357 VDDREF VDDREF pch l=0.26u w=1u
m16045 VDDREF 1360 VDDREF VDDREF pch l=0.26u w=1u
m16046 VDDREF 1361 VDDREF VDDREF pch l=0.26u w=1u
m16047 VDDREF 1363 VDDREF VDDREF pch l=0.26u w=1u
m16048 VDDREF 1366 VDDREF VDDREF pch l=0.26u w=1u
m16049 VDDREF 1367 VDDREF VDDREF pch l=0.26u w=1u
m16050 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m16051 1280 1240 VDDREF VDDREF pch l=0.04u w=0.8u
m16052 1225 1314 VDDREF VDDREF pch l=0.04u w=0.8u
m16053 VDDREF 1346 VDDREF VDDREF pch l=0.26u w=1u
m16054 VDDREF 1347 VDDREF VDDREF pch l=0.26u w=1u
m16055 VDDREF 1350 VDDREF VDDREF pch l=0.26u w=1u
m16056 VDDREF 1351 VDDREF VDDREF pch l=0.26u w=1u
m16057 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16058 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16059 VDDREF 1335 28756 VDDREF pch l=0.04u w=0.24u
m16060 1261 686 VDDREF VDDREF pch l=0.04u w=0.8u
m16061 1262 687 VDDREF VDDREF pch l=0.04u w=0.8u
m16062 VDDREF 1294 1260 VDDREF pch l=0.04u w=0.8u
m16063 VDDREF 417 1267 VDDREF pch l=0.04u w=0.8u
m16064 VDDREF 419 1268 VDDREF pch l=0.04u w=0.8u
m16065 VDDREF 420 1269 VDDREF pch l=0.04u w=0.8u
m16066 VDDREF 422 1270 VDDREF pch l=0.04u w=0.8u
m16067 VDDREF 423 1271 VDDREF pch l=0.04u w=0.8u
m16068 VDDREF 425 1272 VDDREF pch l=0.04u w=0.8u
m16069 1281 1248 VDDREF VDDREF pch l=0.04u w=0.8u
m16070 1282 1249 VDDREF VDDREF pch l=0.04u w=0.8u
m16071 VDDREF 428 1273 VDDREF pch l=0.04u w=0.8u
m16072 VDDREF 429 1274 VDDREF pch l=0.04u w=0.8u
m16073 VDDREF 431 1275 VDDREF pch l=0.04u w=0.8u
m16074 VDDREF 432 1276 VDDREF pch l=0.04u w=0.8u
m16075 VDDREF 433 1277 VDDREF pch l=0.04u w=0.8u
m16076 VDDREF 435 1278 VDDREF pch l=0.04u w=0.8u
m16077 VDDREF 436 1279 VDDREF pch l=0.04u w=0.8u
m16078 VDDREF 683 1280 VDDREF pch l=0.04u w=0.8u
m16079 1266 1313 VDDREF VDDREF pch l=0.04u w=0.8u
m16080 VDDREF 1354 1225 VDDREF pch l=0.04u w=0.8u
m16081 1283 1259 VDDREF VDDREF pch l=0.04u w=0.8u
m16082 28769 1260 VDDREF VDDREF pch l=0.04u w=0.12u
m16083 1267 711 VDDREF VDDREF pch l=0.04u w=0.8u
m16084 1284 1159 VDDREF VDDREF pch l=0.04u w=0.8u
m16085 1268 713 VDDREF VDDREF pch l=0.04u w=0.8u
m16086 1269 714 VDDREF VDDREF pch l=0.04u w=0.8u
m16087 1285 1162 VDDREF VDDREF pch l=0.04u w=0.8u
m16088 1270 716 VDDREF VDDREF pch l=0.04u w=0.8u
m16089 1271 717 VDDREF VDDREF pch l=0.04u w=0.8u
m16090 1286 1165 VDDREF VDDREF pch l=0.04u w=0.8u
m16091 1272 719 VDDREF VDDREF pch l=0.04u w=0.8u
m16092 1287 131 VDDREF VDDREF pch l=0.04u w=0.8u
m16093 1273 722 VDDREF VDDREF pch l=0.04u w=0.8u
m16094 1274 723 VDDREF VDDREF pch l=0.04u w=0.8u
m16095 1288 1169 VDDREF VDDREF pch l=0.04u w=0.8u
m16096 1275 725 VDDREF VDDREF pch l=0.04u w=0.8u
m16097 1276 726 VDDREF VDDREF pch l=0.04u w=0.8u
m16098 1277 727 VDDREF VDDREF pch l=0.04u w=0.8u
m16099 1289 1173 VDDREF VDDREF pch l=0.04u w=0.8u
m16100 1278 729 VDDREF VDDREF pch l=0.04u w=0.8u
m16101 1279 730 VDDREF VDDREF pch l=0.04u w=0.8u
m16102 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16103 VDDREF 1357 VDDREF VDDREF pch l=0.26u w=1u
m16104 VDDREF 1360 VDDREF VDDREF pch l=0.26u w=1u
m16105 VDDREF 1361 VDDREF VDDREF pch l=0.26u w=1u
m16106 VDDREF 1363 VDDREF VDDREF pch l=0.26u w=1u
m16107 VDDREF 1366 VDDREF VDDREF pch l=0.26u w=1u
m16108 VDDREF 1367 VDDREF VDDREF pch l=0.26u w=1u
m16109 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m16110 VDDREF 2648 1266 VDDREF pch l=0.04u w=0.8u
m16111 VDDREF 1346 VDDREF VDDREF pch l=0.26u w=1u
m16112 VDDREF 1347 VDDREF VDDREF pch l=0.26u w=1u
m16113 VDDREF 1350 VDDREF VDDREF pch l=0.26u w=1u
m16114 VDDREF 1351 VDDREF VDDREF pch l=0.26u w=1u
m16115 1225 1354 VDDREF VDDREF pch l=0.04u w=0.8u
m16116 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16117 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16118 1294 1315 28769 VDDREF pch l=0.04u w=0.12u
m16119 1290 1261 VDDREF VDDREF pch l=0.04u w=0.8u
m16120 VDDREF 1190 1284 VDDREF pch l=0.04u w=0.8u
m16121 1291 1262 VDDREF VDDREF pch l=0.04u w=0.8u
m16122 VDDREF 1191 1285 VDDREF pch l=0.04u w=0.8u
m16123 VDDREF 1192 1286 VDDREF pch l=0.04u w=0.8u
m16124 VDDREF 1193 1287 VDDREF pch l=0.04u w=0.8u
m16125 VDDREF 1194 1288 VDDREF pch l=0.04u w=0.8u
m16126 VDDREF 1195 1289 VDDREF pch l=0.04u w=0.8u
m16127 1292 1223 1281 VDDREF pch l=0.04u w=0.8u
m16128 1293 1224 1282 VDDREF pch l=0.04u w=0.8u
m16129 28781 1266 VDDREF VDDREF pch l=0.04u w=0.12u
m16130 1295 1280 VDDREF VDDREF pch l=0.04u w=0.8u
m16131 VDDREF 1314 1225 VDDREF pch l=0.04u w=0.8u
m16132 1296 1372 1294 VDDREF pch l=0.04u w=0.8u
m16133 1297 1110 VDDREF VDDREF pch l=0.04u w=0.8u
m16134 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16135 VDDREF 1357 VDDREF VDDREF pch l=0.26u w=1u
m16136 VDDREF 1360 VDDREF VDDREF pch l=0.26u w=1u
m16137 VDDREF 1361 VDDREF VDDREF pch l=0.26u w=1u
m16138 VDDREF 1363 VDDREF VDDREF pch l=0.26u w=1u
m16139 VDDREF 1366 VDDREF VDDREF pch l=0.26u w=1u
m16140 VDDREF 1367 VDDREF VDDREF pch l=0.26u w=1u
m16141 1298 1267 VDDREF VDDREF pch l=0.04u w=0.8u
m16142 1299 1268 VDDREF VDDREF pch l=0.04u w=0.8u
m16143 1300 1269 VDDREF VDDREF pch l=0.04u w=0.8u
m16144 1301 1270 VDDREF VDDREF pch l=0.04u w=0.8u
m16145 1302 1271 VDDREF VDDREF pch l=0.04u w=0.8u
m16146 1304 1272 VDDREF VDDREF pch l=0.04u w=0.8u
m16147 28786 4328 1292 VDDREF pch l=0.04u w=0.12u
m16148 28787 4328 1293 VDDREF pch l=0.04u w=0.12u
m16149 1305 1273 VDDREF VDDREF pch l=0.04u w=0.8u
m16150 1306 1274 VDDREF VDDREF pch l=0.04u w=0.8u
m16151 1307 1275 VDDREF VDDREF pch l=0.04u w=0.8u
m16152 1308 1276 VDDREF VDDREF pch l=0.04u w=0.8u
m16153 1309 1277 VDDREF VDDREF pch l=0.04u w=0.8u
m16154 1310 1278 VDDREF VDDREF pch l=0.04u w=0.8u
m16155 1311 1279 VDDREF VDDREF pch l=0.04u w=0.8u
m16156 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m16157 1313 1353 28781 VDDREF pch l=0.04u w=0.12u
m16158 VDDREF 1346 VDDREF VDDREF pch l=0.26u w=1u
m16159 VDDREF 1347 VDDREF VDDREF pch l=0.26u w=1u
m16160 VDDREF 1350 VDDREF VDDREF pch l=0.26u w=1u
m16161 VDDREF 1351 VDDREF VDDREF pch l=0.26u w=1u
m16162 1312 1318 1295 VDDREF pch l=0.04u w=0.8u
m16163 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16164 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16165 VDDREF 1283 1297 VDDREF pch l=0.04u w=0.8u
m16166 1316 1290 VDDREF VDDREF pch l=0.04u w=0.8u
m16167 1190 1179 272 VDDREF pch l=0.04u w=0.8u
m16168 1317 1291 VDDREF VDDREF pch l=0.04u w=0.8u
m16169 1191 1184 139 VDDREF pch l=0.04u w=0.8u
m16170 1192 94 FRAC[20] VDDREF pch l=0.04u w=0.8u
m16171 VDDREF 1319 28786 VDDREF pch l=0.04u w=0.12u
m16172 VDDREF 1320 28787 VDDREF pch l=0.04u w=0.12u
m16173 1193 1321 960 VDDREF pch l=0.04u w=0.8u
m16174 1194 960 820 VDDREF pch l=0.04u w=0.8u
m16175 1195 961 FRAC[20] VDDREF pch l=0.04u w=0.8u
m16176 1152 1392 1313 VDDREF pch l=0.04u w=0.8u
m16177 1318 1295 1312 VDDREF pch l=0.04u w=0.8u
m16178 1314 1438 VDDREF VDDREF pch l=0.04u w=0.8u
m16179 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16180 VDDREF 1357 VDDREF VDDREF pch l=0.26u w=1u
m16181 VDDREF 1360 VDDREF VDDREF pch l=0.26u w=1u
m16182 VDDREF 1361 VDDREF VDDREF pch l=0.26u w=1u
m16183 VDDREF 1363 VDDREF VDDREF pch l=0.26u w=1u
m16184 VDDREF 1366 VDDREF VDDREF pch l=0.26u w=1u
m16185 VDDREF 1367 VDDREF VDDREF pch l=0.26u w=1u
m16186 VDDREF 1372 1315 VDDREF pch l=0.04u w=0.8u
m16187 VDDREF 977 1316 VDDREF pch l=0.04u w=0.8u
m16188 1179 272 1190 VDDREF pch l=0.04u w=0.8u
m16189 VDDREF 978 1317 VDDREF pch l=0.04u w=0.8u
m16190 1184 139 1191 VDDREF pch l=0.04u w=0.8u
m16191 94 FRAC[20] 1192 VDDREF pch l=0.04u w=0.8u
m16192 1319 1292 VDDREF VDDREF pch l=0.04u w=0.8u
m16193 1320 1293 VDDREF VDDREF pch l=0.04u w=0.8u
m16194 1321 960 1193 VDDREF pch l=0.04u w=0.8u
m16195 960 820 1194 VDDREF pch l=0.04u w=0.8u
m16196 961 FRAC[20] 1195 VDDREF pch l=0.04u w=0.8u
m16197 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m16198 1322 1298 VDDREF VDDREF pch l=0.04u w=0.8u
m16199 1323 1299 VDDREF VDDREF pch l=0.04u w=0.8u
m16200 1324 1300 VDDREF VDDREF pch l=0.04u w=0.8u
m16201 1325 1301 VDDREF VDDREF pch l=0.04u w=0.8u
m16202 1326 1302 VDDREF VDDREF pch l=0.04u w=0.8u
m16203 1327 1304 VDDREF VDDREF pch l=0.04u w=0.8u
m16204 1328 1305 VDDREF VDDREF pch l=0.04u w=0.8u
m16205 1329 1306 VDDREF VDDREF pch l=0.04u w=0.8u
m16206 1330 1307 VDDREF VDDREF pch l=0.04u w=0.8u
m16207 1331 1308 VDDREF VDDREF pch l=0.04u w=0.8u
m16208 1332 1309 VDDREF VDDREF pch l=0.04u w=0.8u
m16209 1333 1310 VDDREF VDDREF pch l=0.04u w=0.8u
m16210 1334 1311 VDDREF VDDREF pch l=0.04u w=0.8u
m16211 VDDREF 1346 VDDREF VDDREF pch l=0.26u w=1u
m16212 VDDREF 1347 VDDREF VDDREF pch l=0.26u w=1u
m16213 VDDREF 1350 VDDREF VDDREF pch l=0.26u w=1u
m16214 VDDREF 1351 VDDREF VDDREF pch l=0.26u w=1u
m16215 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16216 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16217 VDDREF 1394 1314 VDDREF pch l=0.04u w=0.8u
m16218 1335 1297 VDDREF VDDREF pch l=0.04u w=0.8u
m16219 1316 110 VDDREF VDDREF pch l=0.04u w=0.8u
m16220 1317 293 VDDREF VDDREF pch l=0.04u w=0.8u
m16221 VDDREF 1003 1322 VDDREF pch l=0.04u w=0.8u
m16222 VDDREF 1005 1323 VDDREF pch l=0.04u w=0.8u
m16223 VDDREF 1006 1324 VDDREF pch l=0.04u w=0.8u
m16224 VDDREF 1008 1325 VDDREF pch l=0.04u w=0.8u
m16225 VDDREF 1009 1326 VDDREF pch l=0.04u w=0.8u
m16226 VDDREF 1011 1327 VDDREF pch l=0.04u w=0.8u
m16227 VDDREF 1014 1328 VDDREF pch l=0.04u w=0.8u
m16228 VDDREF 1015 1329 VDDREF pch l=0.04u w=0.8u
m16229 VDDREF 1017 1330 VDDREF pch l=0.04u w=0.8u
m16230 VDDREF 1018 1331 VDDREF pch l=0.04u w=0.8u
m16231 VDDREF 1019 1332 VDDREF pch l=0.04u w=0.8u
m16232 VDDREF 1021 1333 VDDREF pch l=0.04u w=0.8u
m16233 VDDREF 1022 1334 VDDREF pch l=0.04u w=0.8u
m16234 1345 1345 VDDREF VDDREF pch l=0.04u w=1u
m16235 1348 1348 VDDREF VDDREF pch l=0.04u w=1u
m16236 1349 1349 VDDREF VDDREF pch l=0.04u w=1u
m16237 1352 1352 VDDREF VDDREF pch l=0.04u w=1u
m16238 1353 1392 VDDREF VDDREF pch l=0.04u w=0.8u
m16239 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16240 VDDREF 1357 VDDREF VDDREF pch l=0.26u w=1u
m16241 VDDREF 1360 VDDREF VDDREF pch l=0.26u w=1u
m16242 VDDREF 1361 VDDREF VDDREF pch l=0.26u w=1u
m16243 VDDREF 1363 VDDREF VDDREF pch l=0.26u w=1u
m16244 VDDREF 1366 VDDREF VDDREF pch l=0.26u w=1u
m16245 VDDREF 1367 VDDREF VDDREF pch l=0.26u w=1u
m16246 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m16247 VDDREF 1034 1296 VDDREF pch l=0.04u w=0.8u
m16248 1322 21 VDDREF VDDREF pch l=0.04u w=0.8u
m16249 VDDREF 1179 1336 VDDREF pch l=0.04u w=0.8u
m16250 1323 110 VDDREF VDDREF pch l=0.04u w=0.8u
m16251 1324 22 VDDREF VDDREF pch l=0.04u w=0.8u
m16252 VDDREF 1184 1337 VDDREF pch l=0.04u w=0.8u
m16253 1325 313 VDDREF VDDREF pch l=0.04u w=0.8u
m16254 1326 25 VDDREF VDDREF pch l=0.04u w=0.8u
m16255 VDDREF 94 1338 VDDREF pch l=0.04u w=0.8u
m16256 1327 315 VDDREF VDDREF pch l=0.04u w=0.8u
m16257 VDDREF 1319 1339 VDDREF pch l=0.04u w=0.8u
m16258 VDDREF 1320 1340 VDDREF pch l=0.04u w=0.8u
m16259 VDDREF 1321 1341 VDDREF pch l=0.04u w=0.8u
m16260 1328 27 VDDREF VDDREF pch l=0.04u w=0.8u
m16261 1329 28 VDDREF VDDREF pch l=0.04u w=0.8u
m16262 VDDREF 960 1342 VDDREF pch l=0.04u w=0.8u
m16263 1330 131 VDDREF VDDREF pch l=0.04u w=0.8u
m16264 1331 318 VDDREF VDDREF pch l=0.04u w=0.8u
m16265 1332 29 VDDREF VDDREF pch l=0.04u w=0.8u
m16266 VDDREF 961 1343 VDDREF pch l=0.04u w=0.8u
m16267 1333 131 VDDREF VDDREF pch l=0.04u w=0.8u
m16268 1334 318 VDDREF VDDREF pch l=0.04u w=0.8u
m16269 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16270 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16271 1356 377 VDDREF VDDREF pch l=0.04u w=0.8u
m16272 1354 REFDIV[5] VDDREF VDDREF pch l=0.04u w=0.8u
m16273 1358 1358 VDDREF VDDREF pch l=0.04u w=1u
m16274 1359 1359 VDDREF VDDREF pch l=0.04u w=1u
m16275 1362 1362 VDDREF VDDREF pch l=0.04u w=1u
m16276 1364 1364 VDDREF VDDREF pch l=0.04u w=1u
m16277 1365 1365 VDDREF VDDREF pch l=0.04u w=1u
m16278 1368 1368 VDDREF VDDREF pch l=0.04u w=1u
m16279 1369 1511 VDDREF VDDREF pch l=0.04u w=0.8u
m16280 1370 1226 VDDREF VDDREF pch l=0.04u w=0.8u
m16281 1371 1227 VDDREF VDDREF pch l=0.04u w=0.8u
m16282 1001 1339 VDDREF VDDREF pch l=0.04u w=0.8u
m16283 793 1340 VDDREF VDDREF pch l=0.04u w=0.8u
m16284 VDDREF 1392 1355 VDDREF pch l=0.04u w=0.8u
m16285 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16286 VDDREF 377 1354 VDDREF pch l=0.04u w=0.8u
m16287 VDDREF 1395 VDDREF VDDREF pch l=0.26u w=1u
m16288 VDDREF 1372 1369 VDDREF pch l=0.04u w=0.8u
m16289 VDDREF 1316 1370 VDDREF pch l=0.04u w=0.8u
m16290 VDDREF 1317 1371 VDDREF pch l=0.04u w=0.8u
m16291 VDDREF 1404 1372 VDDREF pch l=0.04u w=0.8u
m16292 1379 1242 VDDREF VDDREF pch l=0.04u w=0.8u
m16293 1373 1179 VDDREF VDDREF pch l=0.04u w=0.8u
m16294 1380 1243 VDDREF VDDREF pch l=0.04u w=0.8u
m16295 1381 1244 VDDREF VDDREF pch l=0.04u w=0.8u
m16296 1374 1184 VDDREF VDDREF pch l=0.04u w=0.8u
m16297 1382 1245 VDDREF VDDREF pch l=0.04u w=0.8u
m16298 1383 1246 VDDREF VDDREF pch l=0.04u w=0.8u
m16299 1375 94 VDDREF VDDREF pch l=0.04u w=0.8u
m16300 1384 1247 VDDREF VDDREF pch l=0.04u w=0.8u
m16301 1376 1321 VDDREF VDDREF pch l=0.04u w=0.8u
m16302 1385 1250 VDDREF VDDREF pch l=0.04u w=0.8u
m16303 1386 1251 VDDREF VDDREF pch l=0.04u w=0.8u
m16304 1377 960 VDDREF VDDREF pch l=0.04u w=0.8u
m16305 1387 1252 VDDREF VDDREF pch l=0.04u w=0.8u
m16306 1388 1253 VDDREF VDDREF pch l=0.04u w=0.8u
m16307 1389 1254 VDDREF VDDREF pch l=0.04u w=0.8u
m16308 1378 961 VDDREF VDDREF pch l=0.04u w=0.8u
m16309 1390 1255 VDDREF VDDREF pch l=0.04u w=0.8u
m16310 1391 1256 VDDREF VDDREF pch l=0.04u w=0.8u
m16311 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16312 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16313 1393 377 VDDREF VDDREF pch l=0.04u w=0.8u
m16314 1396 1396 VDDREF VDDREF pch l=0.04u w=1u
m16315 28846 1372 VDDREF VDDREF pch l=0.04u w=0.12u
m16316 VDDREF 1322 1379 VDDREF pch l=0.04u w=0.8u
m16317 VDDREF 272 1373 VDDREF pch l=0.04u w=0.8u
m16318 VDDREF 1323 1380 VDDREF pch l=0.04u w=0.8u
m16319 VDDREF 1324 1381 VDDREF pch l=0.04u w=0.8u
m16320 VDDREF 139 1374 VDDREF pch l=0.04u w=0.8u
m16321 VDDREF 1325 1382 VDDREF pch l=0.04u w=0.8u
m16322 VDDREF 1326 1383 VDDREF pch l=0.04u w=0.8u
m16323 VDDREF FRAC[20] 1375 VDDREF pch l=0.04u w=0.8u
m16324 VDDREF 1327 1384 VDDREF pch l=0.04u w=0.8u
m16325 1397 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16326 1398 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16327 VDDREF 960 1376 VDDREF pch l=0.04u w=0.8u
m16328 VDDREF 1328 1385 VDDREF pch l=0.04u w=0.8u
m16329 VDDREF 1329 1386 VDDREF pch l=0.04u w=0.8u
m16330 VDDREF 820 1377 VDDREF pch l=0.04u w=0.8u
m16331 VDDREF 1330 1387 VDDREF pch l=0.04u w=0.8u
m16332 VDDREF 1331 1388 VDDREF pch l=0.04u w=0.8u
m16333 VDDREF 1332 1389 VDDREF pch l=0.04u w=0.8u
m16334 VDDREF FRAC[20] 1378 VDDREF pch l=0.04u w=0.8u
m16335 VDDREF 1333 1390 VDDREF pch l=0.04u w=0.8u
m16336 VDDREF 1334 1391 VDDREF pch l=0.04u w=0.8u
m16337 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16338 1392 1436 VDDREF VDDREF pch l=0.04u w=0.8u
m16339 VDDREF REFDIV[2] 1393 VDDREF pch l=0.04u w=0.8u
m16340 VDDREF 377 1394 VDDREF pch l=0.04u w=0.8u
m16341 1404 1772 28846 VDDREF pch l=0.04u w=0.12u
m16342 28861 1511 VDDREF VDDREF pch l=0.04u w=0.8u
m16343 VDDREF 1414 VDDREF VDDREF pch l=0.26u w=1u
m16344 VDDREF 1415 VDDREF VDDREF pch l=0.26u w=1u
m16345 1402 346 VDDREF VDDREF pch l=0.04u w=0.8u
m16346 1403 1447 VDDREF VDDREF pch l=0.04u w=0.8u
m16347 VDDREF 2648 1392 VDDREF pch l=0.04u w=0.8u
m16348 VDDREF 1399 1400 VDDREF pch l=0.04u w=1u
m16349 1412 1529 1404 VDDREF pch l=0.04u w=0.8u
m16350 1401 1372 28861 VDDREF pch l=0.04u w=0.8u
m16351 1413 1413 VDDREF VDDREF pch l=0.04u w=1u
m16352 1416 1416 VDDREF VDDREF pch l=0.04u w=1u
m16353 VDDREF 1179 1402 VDDREF pch l=0.04u w=0.8u
m16354 VDDREF 129 1403 VDDREF pch l=0.04u w=0.8u
m16355 VDDREF 1405 1406 VDDREF pch l=0.04u w=1u
m16356 1159 1456 VDDREF VDDREF pch l=0.04u w=0.8u
m16357 1419 1503 VDDREF VDDREF pch l=0.04u w=0.8u
m16358 1162 1457 VDDREF VDDREF pch l=0.04u w=0.8u
m16359 1420 1514 VDDREF VDDREF pch l=0.04u w=0.8u
m16360 1421 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m16361 1422 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m16362 VDDREF 1407 1408 VDDREF pch l=0.04u w=1u
m16363 1423 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m16364 1165 1458 VDDREF VDDREF pch l=0.04u w=0.8u
m16365 1424 FRAC[4] VDDREF VDDREF pch l=0.04u w=0.8u
m16366 1417 4328 1319 VDDREF pch l=0.04u w=0.8u
m16367 1418 4328 1320 VDDREF pch l=0.04u w=0.8u
m16368 VDDREF 1483 1409 VDDREF pch l=0.04u w=0.8u
m16369 1425 1504 VDDREF VDDREF pch l=0.04u w=0.8u
m16370 1426 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16371 1427 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16372 1428 1518 VDDREF VDDREF pch l=0.04u w=0.8u
m16373 1169 1460 VDDREF VDDREF pch l=0.04u w=0.8u
m16374 1429 1519 VDDREF VDDREF pch l=0.04u w=0.8u
m16375 1430 1409 VDDREF VDDREF pch l=0.04u w=0.8u
m16376 1431 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16377 1432 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16378 1433 1522 VDDREF VDDREF pch l=0.04u w=0.8u
m16379 1173 1461 VDDREF VDDREF pch l=0.04u w=0.8u
m16380 1434 FRAC[4] VDDREF VDDREF pch l=0.04u w=0.8u
m16381 1435 1409 VDDREF VDDREF pch l=0.04u w=0.8u
m16382 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16383 1437 1356 VDDREF VDDREF pch l=0.04u w=0.8u
m16384 VDDREF 1411 1410 VDDREF pch l=0.04u w=1u
m16385 VDDREF 1618 1159 VDDREF pch l=0.04u w=0.8u
m16386 VDDREF 1499 1419 VDDREF pch l=0.04u w=0.8u
m16387 VDDREF 1619 1162 VDDREF pch l=0.04u w=0.8u
m16388 VDDREF 1502 1420 VDDREF pch l=0.04u w=0.8u
m16389 VDDREF 1658 1421 VDDREF pch l=0.04u w=0.8u
m16390 VDDREF 1659 1422 VDDREF pch l=0.04u w=0.8u
m16391 VDDREF 1181 1423 VDDREF pch l=0.04u w=0.8u
m16392 VDDREF 1620 1165 VDDREF pch l=0.04u w=0.8u
m16393 VDDREF 1503 1424 VDDREF pch l=0.04u w=0.8u
m16394 28877 1397 1417 VDDREF pch l=0.04u w=0.12u
m16395 28878 1398 1418 VDDREF pch l=0.04u w=0.12u
m16396 VDDREF 131 1425 VDDREF pch l=0.04u w=0.8u
m16397 VDDREF 1504 1428 VDDREF pch l=0.04u w=0.8u
m16398 VDDREF 1621 1169 VDDREF pch l=0.04u w=0.8u
m16399 VDDREF 1505 1429 VDDREF pch l=0.04u w=0.8u
m16400 VDDREF 1506 1430 VDDREF pch l=0.04u w=0.8u
m16401 VDDREF 1507 1433 VDDREF pch l=0.04u w=0.8u
m16402 VDDREF 1622 1173 VDDREF pch l=0.04u w=0.8u
m16403 VDDREF 1508 1434 VDDREF pch l=0.04u w=0.8u
m16404 VDDREF FBDIV[4] 1435 VDDREF pch l=0.04u w=0.8u
m16405 VDDREF 1484 1436 VDDREF pch l=0.04u w=0.8u
m16406 VDDREF 1312 1437 VDDREF pch l=0.04u w=0.8u
m16407 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16408 1438 1463 1090 VDDREF pch l=0.04u w=0.8u
m16409 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16410 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16411 VDDREF 1486 1412 VDDREF pch l=0.04u w=0.8u
m16412 1449 1335 VDDREF VDDREF pch l=0.04u w=0.8u
m16413 VDDREF 1440 1439 VDDREF pch l=0.04u w=1u
m16414 VDDREF 1441 1442 VDDREF pch l=0.04u w=1u
m16415 1450 1179 VDDREF VDDREF pch l=0.04u w=0.8u
m16416 1451 129 VDDREF VDDREF pch l=0.04u w=0.8u
m16417 VDDREF 1466 28877 VDDREF pch l=0.04u w=0.12u
m16418 VDDREF 1467 28878 VDDREF pch l=0.04u w=0.12u
m16419 1459 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16420 1452 4328 1443 VDDREF pch l=0.04u w=0.8u
m16421 1453 4328 1444 VDDREF pch l=0.04u w=0.8u
m16422 1454 4328 1445 VDDREF pch l=0.04u w=0.8u
m16423 1455 4328 1446 VDDREF pch l=0.04u w=0.8u
m16424 VDDREF 1482 VDDREF VDDREF pch l=0.26u w=1u
m16425 VDDREF 2906 1447 VDDREF pch l=0.04u w=0.8u
m16426 28897 1355 VDDREF VDDREF pch l=0.04u w=0.24u
m16427 1463 1090 1438 VDDREF pch l=0.04u w=0.8u
m16428 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16429 28928 1412 VDDREF VDDREF pch l=0.04u w=0.12u
m16430 1466 1417 VDDREF VDDREF pch l=0.04u w=0.8u
m16431 1467 1418 VDDREF VDDREF pch l=0.04u w=0.8u
m16432 VDDREF 2466 1456 VDDREF pch l=0.04u w=0.8u
m16433 1468 1499 VDDREF VDDREF pch l=0.04u w=0.8u
m16434 VDDREF 2468 1457 VDDREF pch l=0.04u w=0.8u
m16435 1469 1502 VDDREF VDDREF pch l=0.04u w=0.8u
m16436 1470 1421 VDDREF VDDREF pch l=0.04u w=0.8u
m16437 1471 1422 VDDREF VDDREF pch l=0.04u w=0.8u
m16438 1472 1423 VDDREF VDDREF pch l=0.04u w=0.8u
m16439 VDDREF 2470 1458 VDDREF pch l=0.04u w=0.8u
m16440 1473 1503 VDDREF VDDREF pch l=0.04u w=0.8u
m16441 1474 131 VDDREF VDDREF pch l=0.04u w=0.8u
m16442 28929 1426 1452 VDDREF pch l=0.04u w=0.12u
m16443 28930 1427 1453 VDDREF pch l=0.04u w=0.12u
m16444 1475 1504 VDDREF VDDREF pch l=0.04u w=0.8u
m16445 VDDREF 2474 1460 VDDREF pch l=0.04u w=0.8u
m16446 1476 1505 VDDREF VDDREF pch l=0.04u w=0.8u
m16447 1477 1506 VDDREF VDDREF pch l=0.04u w=0.8u
m16448 28931 1431 1454 VDDREF pch l=0.04u w=0.12u
m16449 28932 1432 1455 VDDREF pch l=0.04u w=0.12u
m16450 1478 1507 VDDREF VDDREF pch l=0.04u w=0.8u
m16451 VDDREF 2478 1461 VDDREF pch l=0.04u w=0.8u
m16452 1479 1508 VDDREF VDDREF pch l=0.04u w=0.8u
m16453 1480 FBDIV[4] VDDREF VDDREF pch l=0.04u w=0.8u
m16454 1481 1481 VDDREF VDDREF pch l=0.04u w=1u
m16455 1484 1663 28897 VDDREF pch l=0.04u w=0.24u
m16456 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16457 1485 1437 VDDREF VDDREF pch l=0.04u w=0.8u
m16458 VDDREF 1448 1463 VDDREF pch l=0.04u w=0.8u
m16459 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16460 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16461 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16462 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16463 1486 1529 28928 VDDREF pch l=0.04u w=0.12u
m16464 28939 1369 VDDREF VDDREF pch l=0.04u w=0.8u
m16465 1464 346 1179 VDDREF pch l=0.04u w=0.8u
m16466 1456 1671 VDDREF VDDREF pch l=0.04u w=0.8u
m16467 1465 1447 129 VDDREF pch l=0.04u w=0.8u
m16468 1457 1672 VDDREF VDDREF pch l=0.04u w=0.8u
m16469 1458 1673 VDDREF VDDREF pch l=0.04u w=0.8u
m16470 VDDREF 1516 28929 VDDREF pch l=0.04u w=0.12u
m16471 VDDREF 1517 28930 VDDREF pch l=0.04u w=0.12u
m16472 1460 1674 VDDREF VDDREF pch l=0.04u w=0.8u
m16473 VDDREF 1520 28931 VDDREF pch l=0.04u w=0.12u
m16474 VDDREF 1521 28932 VDDREF pch l=0.04u w=0.12u
m16475 1461 1675 VDDREF VDDREF pch l=0.04u w=0.8u
m16476 1491 4328 1483 VDDREF pch l=0.04u w=0.8u
m16477 1510 1623 1484 VDDREF pch l=0.04u w=0.8u
m16478 VDDREF 1393 1485 VDDREF pch l=0.04u w=0.8u
m16479 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16480 1511 1772 1486 VDDREF pch l=0.04u w=0.8u
m16481 1487 1449 28939 VDDREF pch l=0.04u w=0.8u
m16482 346 1179 1464 VDDREF pch l=0.04u w=0.8u
m16483 VDDREF 1531 1456 VDDREF pch l=0.04u w=0.8u
m16484 1447 129 1465 VDDREF pch l=0.04u w=0.8u
m16485 VDDREF 1533 1457 VDDREF pch l=0.04u w=0.8u
m16486 VDDREF 1534 1458 VDDREF pch l=0.04u w=0.8u
m16487 1512 1397 1466 VDDREF pch l=0.04u w=0.8u
m16488 1513 1398 1467 VDDREF pch l=0.04u w=0.8u
m16489 1516 1452 VDDREF VDDREF pch l=0.04u w=0.8u
m16490 1517 1453 VDDREF VDDREF pch l=0.04u w=0.8u
m16491 VDDREF 1535 1460 VDDREF pch l=0.04u w=0.8u
m16492 1520 1454 VDDREF VDDREF pch l=0.04u w=0.8u
m16493 1521 1455 VDDREF VDDREF pch l=0.04u w=0.8u
m16494 VDDREF 1536 1461 VDDREF pch l=0.04u w=0.8u
m16495 1523 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16496 1524 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16497 1525 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16498 1488 1503 1499 VDDREF pch l=0.04u w=0.8u
m16499 VDDREF 1501 1500 VDDREF pch l=0.04u w=1u
m16500 1489 1514 1502 VDDREF pch l=0.04u w=0.8u
m16501 1526 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16502 1527 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16503 1528 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16504 1490 FRAC[4] 1503 VDDREF pch l=0.04u w=0.8u
m16505 28947 1459 1491 VDDREF pch l=0.04u w=0.12u
m16506 1492 1504 131 VDDREF pch l=0.04u w=0.8u
m16507 1493 1518 1504 VDDREF pch l=0.04u w=0.8u
m16508 1494 1519 1505 VDDREF pch l=0.04u w=0.8u
m16509 1495 1409 1506 VDDREF pch l=0.04u w=0.8u
m16510 1496 1522 1507 VDDREF pch l=0.04u w=0.8u
m16511 1497 FRAC[4] 1508 VDDREF pch l=0.04u w=0.8u
m16512 1498 1409 FBDIV[4] VDDREF pch l=0.04u w=0.8u
m16513 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16514 1485 1393 VDDREF VDDREF pch l=0.04u w=0.8u
m16515 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16516 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16517 1448 683 VDDREF VDDREF pch l=0.04u w=0.8u
m16518 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16519 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16520 28956 4328 1512 VDDREF pch l=0.04u w=0.12u
m16521 28957 4328 1513 VDDREF pch l=0.04u w=0.12u
m16522 1503 1499 1488 VDDREF pch l=0.04u w=0.8u
m16523 1514 1502 1489 VDDREF pch l=0.04u w=0.8u
m16524 FRAC[4] 1503 1490 VDDREF pch l=0.04u w=0.8u
m16525 VDDREF 1550 28947 VDDREF pch l=0.04u w=0.12u
m16526 1504 131 1492 VDDREF pch l=0.04u w=0.8u
m16527 1518 1504 1493 VDDREF pch l=0.04u w=0.8u
m16528 1519 1505 1494 VDDREF pch l=0.04u w=0.8u
m16529 1409 1506 1495 VDDREF pch l=0.04u w=0.8u
m16530 1522 1507 1496 VDDREF pch l=0.04u w=0.8u
m16531 FRAC[4] 1508 1497 VDDREF pch l=0.04u w=0.8u
m16532 1409 FBDIV[4] 1498 VDDREF pch l=0.04u w=0.8u
m16533 1510 1572 VDDREF VDDREF pch l=0.04u w=0.8u
m16534 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16535 VDDREF 1437 1485 VDDREF pch l=0.04u w=0.8u
m16536 VDDREF 1561 1448 VDDREF pch l=0.04u w=0.8u
m16537 VDDREF 1772 1529 VDDREF pch l=0.04u w=0.8u
m16538 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16539 VDDREF 1562 28956 VDDREF pch l=0.04u w=0.12u
m16540 VDDREF 1563 28957 VDDREF pch l=0.04u w=0.12u
m16541 1543 1401 VDDREF VDDREF pch l=0.04u w=0.8u
m16542 1530 1464 VDDREF VDDREF pch l=0.04u w=0.8u
m16543 VDDREF 1564 1531 VDDREF pch l=0.04u w=0.8u
m16544 1532 1465 VDDREF VDDREF pch l=0.04u w=0.8u
m16545 VDDREF 1565 1533 VDDREF pch l=0.04u w=0.8u
m16546 VDDREF 1566 1534 VDDREF pch l=0.04u w=0.8u
m16547 1550 1491 VDDREF VDDREF pch l=0.04u w=0.8u
m16548 1539 1426 1516 VDDREF pch l=0.04u w=0.8u
m16549 1540 1427 1517 VDDREF pch l=0.04u w=0.8u
m16550 VDDREF 1567 1535 VDDREF pch l=0.04u w=0.8u
m16551 1541 1431 1520 VDDREF pch l=0.04u w=0.8u
m16552 1542 1432 1521 VDDREF pch l=0.04u w=0.8u
m16553 VDDREF 1568 1536 VDDREF pch l=0.04u w=0.8u
m16554 1544 4328 1537 VDDREF pch l=0.04u w=0.8u
m16555 1545 4328 1538 VDDREF pch l=0.04u w=0.8u
m16556 1546 4328 1180 VDDREF pch l=0.04u w=0.8u
m16557 1547 4328 1470 VDDREF pch l=0.04u w=0.8u
m16558 1548 4328 1471 VDDREF pch l=0.04u w=0.8u
m16559 1549 4328 1472 VDDREF pch l=0.04u w=0.8u
m16560 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16561 VDDREF 2648 1510 VDDREF pch l=0.04u w=0.8u
m16562 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16563 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16564 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16565 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16566 1562 1512 VDDREF VDDREF pch l=0.04u w=0.8u
m16567 1563 1513 VDDREF VDDREF pch l=0.04u w=0.8u
m16568 VDDREF 1335 1543 VDDREF pch l=0.04u w=0.8u
m16569 VDDREF 1370 1530 VDDREF pch l=0.04u w=0.8u
m16570 VDDREF 1371 1532 VDDREF pch l=0.04u w=0.8u
m16571 28968 4328 1539 VDDREF pch l=0.04u w=0.12u
m16572 28969 4328 1540 VDDREF pch l=0.04u w=0.12u
m16573 28970 4328 1541 VDDREF pch l=0.04u w=0.12u
m16574 28971 4328 1542 VDDREF pch l=0.04u w=0.12u
m16575 28972 1523 1544 VDDREF pch l=0.04u w=0.12u
m16576 28973 1524 1545 VDDREF pch l=0.04u w=0.12u
m16577 28974 1525 1546 VDDREF pch l=0.04u w=0.12u
m16578 1551 1488 VDDREF VDDREF pch l=0.04u w=0.8u
m16579 1552 1489 VDDREF VDDREF pch l=0.04u w=0.8u
m16580 28975 1526 1547 VDDREF pch l=0.04u w=0.12u
m16581 28976 1527 1548 VDDREF pch l=0.04u w=0.12u
m16582 28977 1528 1549 VDDREF pch l=0.04u w=0.12u
m16583 1553 1490 VDDREF VDDREF pch l=0.04u w=0.8u
m16584 1554 1492 VDDREF VDDREF pch l=0.04u w=0.8u
m16585 1555 1493 VDDREF VDDREF pch l=0.04u w=0.8u
m16586 1556 1494 VDDREF VDDREF pch l=0.04u w=0.8u
m16587 1557 1495 VDDREF VDDREF pch l=0.04u w=0.8u
m16588 1558 1496 VDDREF VDDREF pch l=0.04u w=0.8u
m16589 1559 1497 VDDREF VDDREF pch l=0.04u w=0.8u
m16590 1560 1498 VDDREF VDDREF pch l=0.04u w=0.8u
m16591 1569 155 VDDREF VDDREF pch l=0.04u w=0.8u
m16592 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16593 28982 1510 VDDREF VDDREF pch l=0.04u w=0.12u
m16594 1570 76 VDDREF VDDREF pch l=0.04u w=0.8u
m16595 VDDREF 1573 1561 VDDREF pch l=0.04u w=0.8u
m16596 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16597 VDDREF 1592 1511 VDDREF pch l=0.04u w=0.8u
m16598 VDDREF 1576 28968 VDDREF pch l=0.04u w=0.12u
m16599 VDDREF 1577 28969 VDDREF pch l=0.04u w=0.12u
m16600 VDDREF 1578 28970 VDDREF pch l=0.04u w=0.12u
m16601 VDDREF 1579 28971 VDDREF pch l=0.04u w=0.12u
m16602 VDDREF 1582 28972 VDDREF pch l=0.04u w=0.12u
m16603 VDDREF 1583 28973 VDDREF pch l=0.04u w=0.12u
m16604 VDDREF 1584 28974 VDDREF pch l=0.04u w=0.12u
m16605 VDDREF 1957 1564 VDDREF pch l=0.04u w=0.8u
m16606 VDDREF 1380 1551 VDDREF pch l=0.04u w=0.8u
m16607 VDDREF 1958 1565 VDDREF pch l=0.04u w=0.8u
m16608 VDDREF 1382 1552 VDDREF pch l=0.04u w=0.8u
m16609 VDDREF 1586 28975 VDDREF pch l=0.04u w=0.12u
m16610 VDDREF 1587 28976 VDDREF pch l=0.04u w=0.12u
m16611 VDDREF 1588 28977 VDDREF pch l=0.04u w=0.12u
m16612 VDDREF 1959 1566 VDDREF pch l=0.04u w=0.8u
m16613 VDDREF 1384 1553 VDDREF pch l=0.04u w=0.8u
m16614 1571 1459 1550 VDDREF pch l=0.04u w=0.8u
m16615 VDDREF 1385 1554 VDDREF pch l=0.04u w=0.8u
m16616 VDDREF 1386 1555 VDDREF pch l=0.04u w=0.8u
m16617 VDDREF 1960 1567 VDDREF pch l=0.04u w=0.8u
m16618 VDDREF 1387 1556 VDDREF pch l=0.04u w=0.8u
m16619 VDDREF 1388 1557 VDDREF pch l=0.04u w=0.8u
m16620 VDDREF 1389 1558 VDDREF pch l=0.04u w=0.8u
m16621 VDDREF 1961 1568 VDDREF pch l=0.04u w=0.8u
m16622 VDDREF 1390 1559 VDDREF pch l=0.04u w=0.8u
m16623 VDDREF 1391 1560 VDDREF pch l=0.04u w=0.8u
m16624 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16625 1572 1623 28982 VDDREF pch l=0.04u w=0.12u
m16626 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16627 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16628 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16629 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16630 28991 1511 VDDREF VDDREF pch l=0.04u w=0.12u
m16631 1574 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16632 1575 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16633 1576 1539 VDDREF VDDREF pch l=0.04u w=0.8u
m16634 1577 1540 VDDREF VDDREF pch l=0.04u w=0.8u
m16635 1578 1541 VDDREF VDDREF pch l=0.04u w=0.8u
m16636 1579 1542 VDDREF VDDREF pch l=0.04u w=0.8u
m16637 1580 1543 VDDREF VDDREF pch l=0.04u w=0.8u
m16638 1581 1530 VDDREF VDDREF pch l=0.04u w=0.8u
m16639 1582 1544 VDDREF VDDREF pch l=0.04u w=0.8u
m16640 1583 1545 VDDREF VDDREF pch l=0.04u w=0.8u
m16641 1584 1546 VDDREF VDDREF pch l=0.04u w=0.8u
m16642 1564 2239 VDDREF VDDREF pch l=0.04u w=0.8u
m16643 1585 1532 VDDREF VDDREF pch l=0.04u w=0.8u
m16644 1565 2240 VDDREF VDDREF pch l=0.04u w=0.8u
m16645 1586 1547 VDDREF VDDREF pch l=0.04u w=0.8u
m16646 1587 1548 VDDREF VDDREF pch l=0.04u w=0.8u
m16647 1588 1549 VDDREF VDDREF pch l=0.04u w=0.8u
m16648 1566 2241 VDDREF VDDREF pch l=0.04u w=0.8u
m16649 28993 4328 1571 VDDREF pch l=0.04u w=0.12u
m16650 1567 2242 VDDREF VDDREF pch l=0.04u w=0.8u
m16651 1568 2243 VDDREF VDDREF pch l=0.04u w=0.8u
m16652 1589 155 VDDREF VDDREF pch l=0.04u w=0.8u
m16653 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16654 1392 1663 1572 VDDREF pch l=0.04u w=0.8u
m16655 1591 76 1485 VDDREF pch l=0.04u w=0.8u
m16656 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16657 VDDREF 1240 1573 VDDREF pch l=0.04u w=0.8u
m16658 1592 1772 28991 VDDREF pch l=0.04u w=0.12u
m16659 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16660 VDDREF 1402 1581 VDDREF pch l=0.04u w=0.8u
m16661 VDDREF 2496 1564 VDDREF pch l=0.04u w=0.8u
m16662 VDDREF 1403 1585 VDDREF pch l=0.04u w=0.8u
m16663 VDDREF 2497 1565 VDDREF pch l=0.04u w=0.8u
m16664 VDDREF 2498 1566 VDDREF pch l=0.04u w=0.8u
m16665 VDDREF 1613 28993 VDDREF pch l=0.04u w=0.12u
m16666 VDDREF 2499 1567 VDDREF pch l=0.04u w=0.8u
m16667 VDDREF 2500 1568 VDDREF pch l=0.04u w=0.8u
m16668 1594 1551 VDDREF VDDREF pch l=0.04u w=0.8u
m16669 1595 1552 VDDREF VDDREF pch l=0.04u w=0.8u
m16670 1596 1553 VDDREF VDDREF pch l=0.04u w=0.8u
m16671 1597 1554 VDDREF VDDREF pch l=0.04u w=0.8u
m16672 1598 1555 VDDREF VDDREF pch l=0.04u w=0.8u
m16673 1599 1556 VDDREF VDDREF pch l=0.04u w=0.8u
m16674 1600 1557 VDDREF VDDREF pch l=0.04u w=0.8u
m16675 1601 1558 VDDREF VDDREF pch l=0.04u w=0.8u
m16676 1602 1559 VDDREF VDDREF pch l=0.04u w=0.8u
m16677 1603 1560 VDDREF VDDREF pch l=0.04u w=0.8u
m16678 VDDREF FBDIV[4] 1589 VDDREF pch l=0.04u w=0.8u
m16679 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16680 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16681 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16682 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16683 29002 1570 1591 VDDREF pch l=0.04u w=0.12u
m16684 1573 2194 VDDREF VDDREF pch l=0.04u w=0.8u
m16685 1604 1696 1592 VDDREF pch l=0.04u w=0.8u
m16686 1605 4328 1562 VDDREF pch l=0.04u w=0.8u
m16687 1606 4328 1563 VDDREF pch l=0.04u w=0.8u
m16688 1613 1571 VDDREF VDDREF pch l=0.04u w=0.8u
m16689 1614 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16690 1615 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16691 1616 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16692 1617 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16693 VDDREF 1637 1593 VDDREF pch l=0.04u w=0.8u
m16694 1607 1523 1582 VDDREF pch l=0.04u w=0.8u
m16695 1608 1524 1583 VDDREF pch l=0.04u w=0.8u
m16696 1609 1525 1584 VDDREF pch l=0.04u w=0.8u
m16697 VDDREF 1419 1594 VDDREF pch l=0.04u w=0.8u
m16698 VDDREF 1420 1595 VDDREF pch l=0.04u w=0.8u
m16699 1610 1526 1586 VDDREF pch l=0.04u w=0.8u
m16700 1611 1527 1587 VDDREF pch l=0.04u w=0.8u
m16701 1612 1528 1588 VDDREF pch l=0.04u w=0.8u
m16702 VDDREF 1424 1596 VDDREF pch l=0.04u w=0.8u
m16703 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16704 VDDREF 1425 1597 VDDREF pch l=0.04u w=0.8u
m16705 VDDREF 1428 1598 VDDREF pch l=0.04u w=0.8u
m16706 VDDREF 1429 1599 VDDREF pch l=0.04u w=0.8u
m16707 VDDREF 1430 1600 VDDREF pch l=0.04u w=0.8u
m16708 VDDREF 1433 1601 VDDREF pch l=0.04u w=0.8u
m16709 VDDREF 1434 1602 VDDREF pch l=0.04u w=0.8u
m16710 VDDREF 1435 1603 VDDREF pch l=0.04u w=0.8u
m16711 1623 1663 VDDREF VDDREF pch l=0.04u w=0.8u
m16712 VDDREF 1631 29002 VDDREF pch l=0.04u w=0.12u
m16713 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16714 VDDREF 1653 1573 VDDREF pch l=0.04u w=0.8u
m16715 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16716 29008 1574 1605 VDDREF pch l=0.04u w=0.12u
m16717 29009 1575 1606 VDDREF pch l=0.04u w=0.12u
m16718 29011 1593 VDDREF VDDREF pch l=0.04u w=0.12u
m16719 1624 1464 VDDREF VDDREF pch l=0.04u w=0.8u
m16720 29012 4328 1607 VDDREF pch l=0.04u w=0.12u
m16721 29013 4328 1608 VDDREF pch l=0.04u w=0.12u
m16722 29014 4328 1609 VDDREF pch l=0.04u w=0.12u
m16723 VDDREF 1719 1618 VDDREF pch l=0.04u w=0.8u
m16724 1625 1465 VDDREF VDDREF pch l=0.04u w=0.8u
m16725 VDDREF 1721 1619 VDDREF pch l=0.04u w=0.8u
m16726 29015 4328 1610 VDDREF pch l=0.04u w=0.12u
m16727 29016 4328 1611 VDDREF pch l=0.04u w=0.12u
m16728 29017 4328 1612 VDDREF pch l=0.04u w=0.12u
m16729 VDDREF 1726 1620 VDDREF pch l=0.04u w=0.8u
m16730 VDDREF 1730 1621 VDDREF pch l=0.04u w=0.8u
m16731 VDDREF 1734 1622 VDDREF pch l=0.04u w=0.8u
m16732 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16733 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16734 1629 1569 VDDREF VDDREF pch l=0.04u w=0.8u
m16735 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16736 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16737 1631 1591 VDDREF VDDREF pch l=0.04u w=0.8u
m16738 VDDREF 1666 1604 VDDREF pch l=0.04u w=0.8u
m16739 VDDREF 1654 29008 VDDREF pch l=0.04u w=0.12u
m16740 VDDREF 1655 29009 VDDREF pch l=0.04u w=0.12u
m16741 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16742 1637 3012 29011 VDDREF pch l=0.04u w=0.12u
m16743 VDDREF 979 29012 VDDREF pch l=0.04u w=0.12u
m16744 VDDREF 1499 29013 VDDREF pch l=0.04u w=0.12u
m16745 VDDREF 1023 29014 VDDREF pch l=0.04u w=0.12u
m16746 VDDREF 1657 29015 VDDREF pch l=0.04u w=0.12u
m16747 VDDREF 1503 29016 VDDREF pch l=0.04u w=0.12u
m16748 VDDREF 1027 29017 VDDREF pch l=0.04u w=0.12u
m16749 1632 4328 1626 VDDREF pch l=0.04u w=0.8u
m16750 1633 4328 1627 VDDREF pch l=0.04u w=0.8u
m16751 1634 4328 1628 VDDREF pch l=0.04u w=0.8u
m16752 1635 4328 1506 VDDREF pch l=0.04u w=0.8u
m16753 1639 1488 VDDREF VDDREF pch l=0.04u w=0.8u
m16754 1641 1489 VDDREF VDDREF pch l=0.04u w=0.8u
m16755 1643 1490 VDDREF VDDREF pch l=0.04u w=0.8u
m16756 1644 1492 VDDREF VDDREF pch l=0.04u w=0.8u
m16757 1645 1493 VDDREF VDDREF pch l=0.04u w=0.8u
m16758 1647 1494 VDDREF VDDREF pch l=0.04u w=0.8u
m16759 1648 1495 VDDREF VDDREF pch l=0.04u w=0.8u
m16760 1649 1496 VDDREF VDDREF pch l=0.04u w=0.8u
m16761 1651 1497 VDDREF VDDREF pch l=0.04u w=0.8u
m16762 1652 1498 VDDREF VDDREF pch l=0.04u w=0.8u
m16763 VDDREF 1613 1629 VDDREF pch l=0.04u w=0.8u
m16764 VDDREF 1663 1630 VDDREF pch l=0.04u w=0.8u
m16765 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16766 1653 1677 VDDREF VDDREF pch l=0.04u w=0.8u
m16767 VDDREF 1664 VDDREF VDDREF pch l=0.26u w=1u
m16768 29029 1604 VDDREF VDDREF pch l=0.04u w=0.12u
m16769 1654 1605 VDDREF VDDREF pch l=0.04u w=0.8u
m16770 1655 1606 VDDREF VDDREF pch l=0.04u w=0.8u
m16771 1656 1744 1637 VDDREF pch l=0.04u w=0.8u
m16772 979 1607 VDDREF VDDREF pch l=0.04u w=0.8u
m16773 1499 1608 VDDREF VDDREF pch l=0.04u w=0.8u
m16774 VDDREF 1667 VDDREF VDDREF pch l=0.26u w=1u
m16775 1023 1609 VDDREF VDDREF pch l=0.04u w=0.8u
m16776 1657 1610 VDDREF VDDREF pch l=0.04u w=0.8u
m16777 1503 1611 VDDREF VDDREF pch l=0.04u w=0.8u
m16778 VDDREF 1669 VDDREF VDDREF pch l=0.26u w=1u
m16779 1027 1612 VDDREF VDDREF pch l=0.04u w=0.8u
m16780 29032 1614 1632 VDDREF pch l=0.04u w=0.12u
m16781 29033 1615 1633 VDDREF pch l=0.04u w=0.12u
m16782 29034 1616 1634 VDDREF pch l=0.04u w=0.12u
m16783 29035 1617 1635 VDDREF pch l=0.04u w=0.12u
m16784 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16785 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16786 1636 1370 1464 VDDREF pch l=0.04u w=0.8u
m16787 1537 1671 1638 VDDREF pch l=0.04u w=0.8u
m16788 138 1371 1465 VDDREF pch l=0.04u w=0.8u
m16789 1658 1672 1640 VDDREF pch l=0.04u w=0.8u
m16790 1660 1673 1642 VDDREF pch l=0.04u w=0.8u
m16791 1444 1674 1646 VDDREF pch l=0.04u w=0.8u
m16792 1446 1675 1650 VDDREF pch l=0.04u w=0.8u
m16793 1662 1570 1631 VDDREF pch l=0.04u w=0.8u
m16794 VDDREF 1677 1653 VDDREF pch l=0.04u w=0.8u
m16795 1665 1665 VDDREF VDDREF pch l=0.04u w=1u
m16796 VDDREF 1681 VDDREF VDDREF pch l=0.26u w=1u
m16797 1666 1696 29029 VDDREF pch l=0.04u w=0.12u
m16798 1668 1668 VDDREF VDDREF pch l=0.04u w=1u
m16799 1670 1670 VDDREF VDDREF pch l=0.04u w=1u
m16800 VDDREF 1685 29032 VDDREF pch l=0.04u w=0.12u
m16801 VDDREF 1686 29033 VDDREF pch l=0.04u w=0.12u
m16802 VDDREF 1687 29034 VDDREF pch l=0.04u w=0.12u
m16803 VDDREF 1688 29035 VDDREF pch l=0.04u w=0.12u
m16804 1370 1464 1636 VDDREF pch l=0.04u w=0.8u
m16805 1671 1638 1537 VDDREF pch l=0.04u w=0.8u
m16806 1371 1465 138 VDDREF pch l=0.04u w=0.8u
m16807 1672 1640 1658 VDDREF pch l=0.04u w=0.8u
m16808 1673 1642 1660 VDDREF pch l=0.04u w=0.8u
m16809 1674 1646 1444 VDDREF pch l=0.04u w=0.8u
m16810 1675 1650 1446 VDDREF pch l=0.04u w=0.8u
m16811 1538 1380 1488 VDDREF pch l=0.04u w=0.8u
m16812 1659 1382 1489 VDDREF pch l=0.04u w=0.8u
m16813 1502 1384 1490 VDDREF pch l=0.04u w=0.8u
m16814 1483 1385 1492 VDDREF pch l=0.04u w=0.8u
m16815 1627 1386 1493 VDDREF pch l=0.04u w=0.8u
m16816 1661 1387 1494 VDDREF pch l=0.04u w=0.8u
m16817 1518 1388 1495 VDDREF pch l=0.04u w=0.8u
m16818 1506 1389 1496 VDDREF pch l=0.04u w=0.8u
m16819 1519 1390 1497 VDDREF pch l=0.04u w=0.8u
m16820 1522 1391 1498 VDDREF pch l=0.04u w=0.8u
m16821 1676 1629 VDDREF VDDREF pch l=0.04u w=0.8u
m16822 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16823 1663 1708 VDDREF VDDREF pch l=0.04u w=0.8u
m16824 29051 76 1662 VDDREF pch l=0.04u w=0.12u
m16825 1680 1680 VDDREF VDDREF pch l=0.04u w=1u
m16826 1682 1772 1666 VDDREF pch l=0.04u w=0.8u
m16827 VDDREF 1698 VDDREF VDDREF pch l=0.26u w=1u
m16828 VDDREF 1699 VDDREF VDDREF pch l=0.26u w=1u
m16829 1683 1574 1654 VDDREF pch l=0.04u w=0.8u
m16830 1684 1575 1655 VDDREF pch l=0.04u w=0.8u
m16831 1685 1632 VDDREF VDDREF pch l=0.04u w=0.8u
m16832 1686 1633 VDDREF VDDREF pch l=0.04u w=0.8u
m16833 1687 1634 VDDREF VDDREF pch l=0.04u w=0.8u
m16834 1688 1635 VDDREF VDDREF pch l=0.04u w=0.8u
m16835 VDDREF 1718 1656 VDDREF pch l=0.04u w=0.8u
m16836 1380 1488 1538 VDDREF pch l=0.04u w=0.8u
m16837 1382 1489 1659 VDDREF pch l=0.04u w=0.8u
m16838 1384 1490 1502 VDDREF pch l=0.04u w=0.8u
m16839 1385 1492 1483 VDDREF pch l=0.04u w=0.8u
m16840 1386 1493 1627 VDDREF pch l=0.04u w=0.8u
m16841 1387 1494 1661 VDDREF pch l=0.04u w=0.8u
m16842 1388 1495 1518 VDDREF pch l=0.04u w=0.8u
m16843 1389 1496 1506 VDDREF pch l=0.04u w=0.8u
m16844 1390 1497 1519 VDDREF pch l=0.04u w=0.8u
m16845 1391 1498 1522 VDDREF pch l=0.04u w=0.8u
m16846 VDDREF 1589 1676 VDDREF pch l=0.04u w=0.8u
m16847 VDDREF 2648 1663 VDDREF pch l=0.04u w=0.8u
m16848 VDDREF 1318 29051 VDDREF pch l=0.04u w=0.12u
m16849 VDDREF 1737 1677 VDDREF pch l=0.04u w=0.8u
m16850 VDDREF 1678 1679 VDDREF pch l=0.04u w=1u
m16851 1697 1697 VDDREF VDDREF pch l=0.04u w=1u
m16852 1700 1700 VDDREF VDDREF pch l=0.04u w=1u
m16853 29066 4328 1683 VDDREF pch l=0.04u w=0.12u
m16854 29067 4328 1684 VDDREF pch l=0.04u w=0.12u
m16855 29070 1656 VDDREF VDDREF pch l=0.04u w=0.12u
m16856 1701 110 VDDREF VDDREF pch l=0.04u w=0.8u
m16857 VDDREF 1671 1689 VDDREF pch l=0.04u w=0.8u
m16858 1702 1741 VDDREF VDDREF pch l=0.04u w=0.8u
m16859 VDDREF 1672 1690 VDDREF pch l=0.04u w=0.8u
m16860 VDDREF 1673 1691 VDDREF pch l=0.04u w=0.8u
m16861 VDDREF 1674 1692 VDDREF pch l=0.04u w=0.8u
m16862 VDDREF 1675 1693 VDDREF pch l=0.04u w=0.8u
m16863 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16864 1318 1662 VDDREF VDDREF pch l=0.04u w=0.8u
m16865 29076 1677 VDDREF VDDREF pch l=0.04u w=0.12u
m16866 VDDREF 1695 1694 VDDREF pch l=0.04u w=1u
m16867 VDDREF 1772 1696 VDDREF pch l=0.04u w=0.8u
m16868 VDDREF 1738 29066 VDDREF pch l=0.04u w=0.12u
m16869 VDDREF 1739 29067 VDDREF pch l=0.04u w=0.12u
m16870 1718 1744 29070 VDDREF pch l=0.04u w=0.12u
m16871 1710 1614 1685 VDDREF pch l=0.04u w=0.8u
m16872 1711 1615 1686 VDDREF pch l=0.04u w=0.8u
m16873 1712 1616 1687 VDDREF pch l=0.04u w=0.8u
m16874 1713 1617 1688 VDDREF pch l=0.04u w=0.8u
m16875 VDDREF 888 1701 VDDREF pch l=0.04u w=0.8u
m16876 VDDREF 441 1702 VDDREF pch l=0.04u w=0.8u
m16877 VDDREF 1703 1704 VDDREF pch l=0.04u w=1u
m16878 1720 1791 VDDREF VDDREF pch l=0.04u w=0.8u
m16879 1722 1803 VDDREF VDDREF pch l=0.04u w=0.8u
m16880 1723 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m16881 1724 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m16882 VDDREF 1705 1706 VDDREF pch l=0.04u w=1u
m16883 1725 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m16884 1727 FRAC[5] VDDREF VDDREF pch l=0.04u w=0.8u
m16885 VDDREF 1770 1707 VDDREF pch l=0.04u w=0.8u
m16886 1728 1792 VDDREF VDDREF pch l=0.04u w=0.8u
m16887 1729 1805 VDDREF VDDREF pch l=0.04u w=0.8u
m16888 1731 1628 VDDREF VDDREF pch l=0.04u w=0.8u
m16889 1732 1707 VDDREF VDDREF pch l=0.04u w=0.8u
m16890 1733 1806 VDDREF VDDREF pch l=0.04u w=0.8u
m16891 1735 FRAC[5] VDDREF VDDREF pch l=0.04u w=0.8u
m16892 1736 1707 VDDREF VDDREF pch l=0.04u w=0.8u
m16893 VDDREF 1750 1708 VDDREF pch l=0.04u w=0.8u
m16894 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m16895 1737 76 29076 VDDREF pch l=0.04u w=0.12u
m16896 1738 1683 VDDREF VDDREF pch l=0.04u w=0.8u
m16897 1739 1684 VDDREF VDDREF pch l=0.04u w=0.8u
m16898 1740 3012 1718 VDDREF pch l=0.04u w=0.8u
m16899 VDDREF 1715 1714 VDDREF pch l=0.04u w=1u
m16900 VDDREF 1716 1717 VDDREF pch l=0.04u w=1u
m16901 29089 4328 1710 VDDREF pch l=0.04u w=0.12u
m16902 29090 4328 1711 VDDREF pch l=0.04u w=0.12u
m16903 29091 4328 1712 VDDREF pch l=0.04u w=0.12u
m16904 29092 4328 1713 VDDREF pch l=0.04u w=0.12u
m16905 VDDREF 1746 VDDREF VDDREF pch l=0.26u w=1u
m16906 1719 1879 VDDREF VDDREF pch l=0.04u w=0.8u
m16907 VDDREF 1789 1720 VDDREF pch l=0.04u w=0.8u
m16908 1721 1881 VDDREF VDDREF pch l=0.04u w=0.8u
m16909 VDDREF 1790 1722 VDDREF pch l=0.04u w=0.8u
m16910 VDDREF 1944 1723 VDDREF pch l=0.04u w=0.8u
m16911 VDDREF 1945 1724 VDDREF pch l=0.04u w=0.8u
m16912 VDDREF 892 1725 VDDREF pch l=0.04u w=0.8u
m16913 1726 1883 VDDREF VDDREF pch l=0.04u w=0.8u
m16914 VDDREF 1791 1727 VDDREF pch l=0.04u w=0.8u
m16915 VDDREF 131 1728 VDDREF pch l=0.04u w=0.8u
m16916 VDDREF 1792 1729 VDDREF pch l=0.04u w=0.8u
m16917 1730 1887 VDDREF VDDREF pch l=0.04u w=0.8u
m16918 VDDREF 1753 1731 VDDREF pch l=0.04u w=0.8u
m16919 VDDREF 1793 1732 VDDREF pch l=0.04u w=0.8u
m16920 VDDREF 1794 1733 VDDREF pch l=0.04u w=0.8u
m16921 1734 1891 VDDREF VDDREF pch l=0.04u w=0.8u
m16922 VDDREF 1754 1735 VDDREF pch l=0.04u w=0.8u
m16923 VDDREF FBDIV[5] 1736 VDDREF pch l=0.04u w=0.8u
m16924 29093 1630 VDDREF VDDREF pch l=0.04u w=0.24u
m16925 1742 1318 VDDREF VDDREF pch l=0.04u w=0.8u
m16926 1743 1844 1737 VDDREF pch l=0.04u w=0.8u
m16927 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m16928 VDDREF 1372 1682 VDDREF pch l=0.04u w=0.8u
m16929 VDDREF 1753 29089 VDDREF pch l=0.04u w=0.12u
m16930 VDDREF 1504 29090 VDDREF pch l=0.04u w=0.12u
m16931 VDDREF 1754 29091 VDDREF pch l=0.04u w=0.12u
m16932 VDDREF 1507 29092 VDDREF pch l=0.04u w=0.12u
m16933 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m16934 1745 1745 VDDREF VDDREF pch l=0.04u w=1u
m16935 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m16936 1747 888 VDDREF VDDREF pch l=0.04u w=0.8u
m16937 VDDREF 1773 1719 VDDREF pch l=0.04u w=0.8u
m16938 1748 441 VDDREF VDDREF pch l=0.04u w=0.8u
m16939 VDDREF 1775 1721 VDDREF pch l=0.04u w=0.8u
m16940 VDDREF 1777 1726 VDDREF pch l=0.04u w=0.8u
m16941 VDDREF 1782 1730 VDDREF pch l=0.04u w=0.8u
m16942 VDDREF 1786 1734 VDDREF pch l=0.04u w=0.8u
m16943 1749 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16944 VDDREF 3180 1741 VDDREF pch l=0.04u w=0.8u
m16945 1750 1934 29093 VDDREF pch l=0.04u w=0.24u
m16946 VDDREF 1318 1742 VDDREF pch l=0.04u w=0.8u
m16947 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m16948 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m16949 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m16950 1751 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16951 1752 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16952 1753 1710 VDDREF VDDREF pch l=0.04u w=0.8u
m16953 1504 1711 VDDREF VDDREF pch l=0.04u w=0.8u
m16954 1754 1712 VDDREF VDDREF pch l=0.04u w=0.8u
m16955 1507 1713 VDDREF VDDREF pch l=0.04u w=0.8u
m16956 VDDREF 3012 1744 VDDREF pch l=0.04u w=0.8u
m16957 1757 1789 VDDREF VDDREF pch l=0.04u w=0.8u
m16958 1758 1790 VDDREF VDDREF pch l=0.04u w=0.8u
m16959 1759 1723 VDDREF VDDREF pch l=0.04u w=0.8u
m16960 1760 1724 VDDREF VDDREF pch l=0.04u w=0.8u
m16961 1761 1725 VDDREF VDDREF pch l=0.04u w=0.8u
m16962 1762 1791 VDDREF VDDREF pch l=0.04u w=0.8u
m16963 1763 131 VDDREF VDDREF pch l=0.04u w=0.8u
m16964 1764 1792 VDDREF VDDREF pch l=0.04u w=0.8u
m16965 1765 1753 VDDREF VDDREF pch l=0.04u w=0.8u
m16966 1766 1793 VDDREF VDDREF pch l=0.04u w=0.8u
m16967 1767 1794 VDDREF VDDREF pch l=0.04u w=0.8u
m16968 1768 1754 VDDREF VDDREF pch l=0.04u w=0.8u
m16969 1769 FBDIV[5] VDDREF VDDREF pch l=0.04u w=0.8u
m16970 1771 1894 1750 VDDREF pch l=0.04u w=0.8u
m16971 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m16972 VDDREF 1813 1743 VDDREF pch l=0.04u w=0.8u
m16973 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m16974 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m16975 1772 1848 VDDREF VDDREF pch l=0.04u w=0.8u
m16976 1755 110 888 VDDREF pch l=0.04u w=0.8u
m16977 1773 1638 VDDREF VDDREF pch l=0.04u w=0.8u
m16978 1756 1741 441 VDDREF pch l=0.04u w=0.8u
m16979 1775 1640 VDDREF VDDREF pch l=0.04u w=0.8u
m16980 1777 1642 VDDREF VDDREF pch l=0.04u w=0.8u
m16981 1782 1646 VDDREF VDDREF pch l=0.04u w=0.8u
m16982 1786 1650 VDDREF VDDREF pch l=0.04u w=0.8u
m16983 1779 4328 1770 VDDREF pch l=0.04u w=0.8u
m16984 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m16985 1796 1742 VDDREF VDDREF pch l=0.04u w=0.8u
m16986 29119 1743 VDDREF VDDREF pch l=0.04u w=0.12u
m16987 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m16988 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m16989 VDDREF 1848 1772 VDDREF pch l=0.04u w=0.8u
m16990 1797 4328 1738 VDDREF pch l=0.04u w=0.8u
m16991 1798 4328 1739 VDDREF pch l=0.04u w=0.8u
m16992 1799 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16993 1800 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16994 1801 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16995 1802 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m16996 VDDREF 1826 1740 VDDREF pch l=0.04u w=0.8u
m16997 110 888 1755 VDDREF pch l=0.04u w=0.8u
m16998 VDDREF 1671 1773 VDDREF pch l=0.04u w=0.8u
m16999 1741 441 1756 VDDREF pch l=0.04u w=0.8u
m17000 VDDREF 1672 1775 VDDREF pch l=0.04u w=0.8u
m17001 VDDREF 1673 1777 VDDREF pch l=0.04u w=0.8u
m17002 VDDREF 1674 1782 VDDREF pch l=0.04u w=0.8u
m17003 VDDREF 1675 1786 VDDREF pch l=0.04u w=0.8u
m17004 1807 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17005 1808 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17006 1809 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17007 1774 1791 1789 VDDREF pch l=0.04u w=0.8u
m17008 1776 1803 1790 VDDREF pch l=0.04u w=0.8u
m17009 1810 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17010 1811 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17011 1812 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17012 1778 FRAC[5] 1791 VDDREF pch l=0.04u w=0.8u
m17013 29126 1749 1779 VDDREF pch l=0.04u w=0.12u
m17014 1780 1792 131 VDDREF pch l=0.04u w=0.8u
m17015 1781 1805 1792 VDDREF pch l=0.04u w=0.8u
m17016 1783 1628 1753 VDDREF pch l=0.04u w=0.8u
m17017 1784 1707 1793 VDDREF pch l=0.04u w=0.8u
m17018 1785 1806 1794 VDDREF pch l=0.04u w=0.8u
m17019 1787 FRAC[5] 1754 VDDREF pch l=0.04u w=0.8u
m17020 1788 1707 FBDIV[5] VDDREF pch l=0.04u w=0.8u
m17021 1771 1851 VDDREF VDDREF pch l=0.04u w=0.8u
m17022 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m17023 VDDREF 1240 1796 VDDREF pch l=0.04u w=0.8u
m17024 1813 1844 29119 VDDREF pch l=0.04u w=0.12u
m17025 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m17026 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m17027 1772 1848 VDDREF VDDREF pch l=0.04u w=0.8u
m17028 29131 1751 1797 VDDREF pch l=0.04u w=0.12u
m17029 29132 1752 1798 VDDREF pch l=0.04u w=0.12u
m17030 29133 1740 VDDREF VDDREF pch l=0.04u w=0.12u
m17031 1791 1789 1774 VDDREF pch l=0.04u w=0.8u
m17032 1803 1790 1776 VDDREF pch l=0.04u w=0.8u
m17033 FRAC[5] 1791 1778 VDDREF pch l=0.04u w=0.8u
m17034 VDDREF 1833 29126 VDDREF pch l=0.04u w=0.12u
m17035 1792 131 1780 VDDREF pch l=0.04u w=0.8u
m17036 1805 1792 1781 VDDREF pch l=0.04u w=0.8u
m17037 1628 1753 1783 VDDREF pch l=0.04u w=0.8u
m17038 1707 1793 1784 VDDREF pch l=0.04u w=0.8u
m17039 1806 1794 1785 VDDREF pch l=0.04u w=0.8u
m17040 FRAC[5] 1754 1787 VDDREF pch l=0.04u w=0.8u
m17041 1707 FBDIV[5] 1788 VDDREF pch l=0.04u w=0.8u
m17042 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m17043 VDDREF 2648 1771 VDDREF pch l=0.04u w=0.8u
m17044 1796 683 VDDREF VDDREF pch l=0.04u w=0.8u
m17045 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m17046 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m17047 1821 76 1813 VDDREF pch l=0.04u w=0.8u
m17048 VDDREF 1848 1772 VDDREF pch l=0.04u w=0.8u
m17049 VDDREF 1846 29131 VDDREF pch l=0.04u w=0.12u
m17050 VDDREF 1847 29132 VDDREF pch l=0.04u w=0.12u
m17051 1826 3012 29133 VDDREF pch l=0.04u w=0.12u
m17052 1822 4328 1814 VDDREF pch l=0.04u w=0.8u
m17053 1823 4328 1661 VDDREF pch l=0.04u w=0.8u
m17054 1824 4328 1815 VDDREF pch l=0.04u w=0.8u
m17055 1825 4328 1519 VDDREF pch l=0.04u w=0.8u
m17056 1816 1755 VDDREF VDDREF pch l=0.04u w=0.8u
m17057 1671 979 1657 VDDREF pch l=0.04u w=0.8u
m17058 1817 1756 VDDREF VDDREF pch l=0.04u w=0.8u
m17059 1672 1660 139 VDDREF pch l=0.04u w=0.8u
m17060 1673 1657 FRAC[19] VDDREF pch l=0.04u w=0.8u
m17061 1833 1779 VDDREF VDDREF pch l=0.04u w=0.8u
m17062 1674 1577 1446 VDDREF pch l=0.04u w=0.8u
m17063 1675 1579 FRAC[19] VDDREF pch l=0.04u w=0.8u
m17064 1827 4328 1819 VDDREF pch l=0.04u w=0.8u
m17065 1828 4328 1820 VDDREF pch l=0.04u w=0.8u
m17066 1829 4328 891 VDDREF pch l=0.04u w=0.8u
m17067 1830 4328 1759 VDDREF pch l=0.04u w=0.8u
m17068 1831 4328 1760 VDDREF pch l=0.04u w=0.8u
m17069 1832 4328 1761 VDDREF pch l=0.04u w=0.8u
m17070 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m17071 29142 1771 VDDREF VDDREF pch l=0.04u w=0.12u
m17072 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m17073 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m17074 1846 1797 VDDREF VDDREF pch l=0.04u w=0.8u
m17075 1847 1798 VDDREF VDDREF pch l=0.04u w=0.8u
m17076 1849 1917 1826 VDDREF pch l=0.04u w=0.8u
m17077 29148 1799 1822 VDDREF pch l=0.04u w=0.12u
m17078 29149 1800 1823 VDDREF pch l=0.04u w=0.12u
m17079 29150 1801 1824 VDDREF pch l=0.04u w=0.12u
m17080 29151 1802 1825 VDDREF pch l=0.04u w=0.12u
m17081 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m17082 VDDREF 1581 1816 VDDREF pch l=0.04u w=0.8u
m17083 979 1657 1671 VDDREF pch l=0.04u w=0.8u
m17084 VDDREF 1585 1817 VDDREF pch l=0.04u w=0.8u
m17085 1660 139 1672 VDDREF pch l=0.04u w=0.8u
m17086 1657 FRAC[19] 1673 VDDREF pch l=0.04u w=0.8u
m17087 1577 1446 1674 VDDREF pch l=0.04u w=0.8u
m17088 1579 FRAC[19] 1675 VDDREF pch l=0.04u w=0.8u
m17089 29152 1807 1827 VDDREF pch l=0.04u w=0.12u
m17090 29153 1808 1828 VDDREF pch l=0.04u w=0.12u
m17091 29154 1809 1829 VDDREF pch l=0.04u w=0.12u
m17092 1834 1774 VDDREF VDDREF pch l=0.04u w=0.8u
m17093 1835 1776 VDDREF VDDREF pch l=0.04u w=0.8u
m17094 29155 1810 1830 VDDREF pch l=0.04u w=0.12u
m17095 29156 1811 1831 VDDREF pch l=0.04u w=0.12u
m17096 29157 1812 1832 VDDREF pch l=0.04u w=0.12u
m17097 1836 1778 VDDREF VDDREF pch l=0.04u w=0.8u
m17098 1837 1780 VDDREF VDDREF pch l=0.04u w=0.8u
m17099 1838 1781 VDDREF VDDREF pch l=0.04u w=0.8u
m17100 1839 1783 VDDREF VDDREF pch l=0.04u w=0.8u
m17101 1840 1784 VDDREF VDDREF pch l=0.04u w=0.8u
m17102 1841 1785 VDDREF VDDREF pch l=0.04u w=0.8u
m17103 1842 1787 VDDREF VDDREF pch l=0.04u w=0.8u
m17104 1843 1788 VDDREF VDDREF pch l=0.04u w=0.8u
m17105 1850 155 VDDREF VDDREF pch l=0.04u w=0.8u
m17106 1851 1894 29142 VDDREF pch l=0.04u w=0.12u
m17107 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m17108 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m17109 1852 1796 VDDREF VDDREF pch l=0.04u w=0.8u
m17110 1853 1943 VDDREF VDDREF pch l=0.04u w=0.8u
m17111 VDDREF 76 1844 VDDREF pch l=0.04u w=0.8u
m17112 1848 1916 VDDREF VDDREF pch l=0.04u w=0.8u
m17113 VDDREF 1863 29148 VDDREF pch l=0.04u w=0.12u
m17114 VDDREF 1864 29149 VDDREF pch l=0.04u w=0.12u
m17115 VDDREF 1865 29150 VDDREF pch l=0.04u w=0.12u
m17116 VDDREF 1866 29151 VDDREF pch l=0.04u w=0.12u
m17117 VDDREF 1868 29152 VDDREF pch l=0.04u w=0.12u
m17118 VDDREF 1869 29153 VDDREF pch l=0.04u w=0.12u
m17119 VDDREF 1870 29154 VDDREF pch l=0.04u w=0.12u
m17120 VDDREF 1594 1834 VDDREF pch l=0.04u w=0.8u
m17121 VDDREF 1595 1835 VDDREF pch l=0.04u w=0.8u
m17122 VDDREF 1872 29155 VDDREF pch l=0.04u w=0.12u
m17123 VDDREF 1873 29156 VDDREF pch l=0.04u w=0.12u
m17124 VDDREF 1874 29157 VDDREF pch l=0.04u w=0.12u
m17125 VDDREF 1596 1836 VDDREF pch l=0.04u w=0.8u
m17126 1854 1749 1833 VDDREF pch l=0.04u w=0.8u
m17127 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m17128 VDDREF 1597 1837 VDDREF pch l=0.04u w=0.8u
m17129 VDDREF 1598 1838 VDDREF pch l=0.04u w=0.8u
m17130 VDDREF 1599 1839 VDDREF pch l=0.04u w=0.8u
m17131 VDDREF 1600 1840 VDDREF pch l=0.04u w=0.8u
m17132 VDDREF 1601 1841 VDDREF pch l=0.04u w=0.8u
m17133 VDDREF 1602 1842 VDDREF pch l=0.04u w=0.8u
m17134 VDDREF 1603 1843 VDDREF pch l=0.04u w=0.8u
m17135 1663 1934 1851 VDDREF pch l=0.04u w=0.8u
m17136 1860 1876 1852 VDDREF pch l=0.04u w=0.8u
m17137 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m17138 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m17139 VDDREF 1878 1848 VDDREF pch l=0.04u w=0.8u
m17140 1861 1751 1846 VDDREF pch l=0.04u w=0.8u
m17141 1862 1752 1847 VDDREF pch l=0.04u w=0.8u
m17142 1863 1822 VDDREF VDDREF pch l=0.04u w=0.8u
m17143 1864 1823 VDDREF VDDREF pch l=0.04u w=0.8u
m17144 1865 1824 VDDREF VDDREF pch l=0.04u w=0.8u
m17145 1866 1825 VDDREF VDDREF pch l=0.04u w=0.8u
m17146 VDDREF 1899 1849 VDDREF pch l=0.04u w=0.8u
m17147 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m17148 1867 1816 VDDREF VDDREF pch l=0.04u w=0.8u
m17149 1868 1827 VDDREF VDDREF pch l=0.04u w=0.8u
m17150 1869 1828 VDDREF VDDREF pch l=0.04u w=0.8u
m17151 1870 1829 VDDREF VDDREF pch l=0.04u w=0.8u
m17152 VDDREF 979 1855 VDDREF pch l=0.04u w=0.8u
m17153 1871 1817 VDDREF VDDREF pch l=0.04u w=0.8u
m17154 VDDREF 1660 1856 VDDREF pch l=0.04u w=0.8u
m17155 1872 1830 VDDREF VDDREF pch l=0.04u w=0.8u
m17156 1873 1831 VDDREF VDDREF pch l=0.04u w=0.8u
m17157 1874 1832 VDDREF VDDREF pch l=0.04u w=0.8u
m17158 VDDREF 1657 1857 VDDREF pch l=0.04u w=0.8u
m17159 29167 4328 1854 VDDREF pch l=0.04u w=0.12u
m17160 VDDREF 1577 1858 VDDREF pch l=0.04u w=0.8u
m17161 VDDREF 1579 1859 VDDREF pch l=0.04u w=0.8u
m17162 1875 155 VDDREF VDDREF pch l=0.04u w=0.8u
m17163 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m17164 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m17165 1876 1852 1860 VDDREF pch l=0.04u w=0.8u
m17166 1877 1657 VDDREF VDDREF pch l=0.04u w=0.8u
m17167 1821 1936 VDDREF VDDREF pch l=0.04u w=0.8u
m17168 29173 4328 1861 VDDREF pch l=0.04u w=0.12u
m17169 29174 4328 1862 VDDREF pch l=0.04u w=0.12u
m17170 29176 1849 VDDREF VDDREF pch l=0.04u w=0.12u
m17171 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m17172 VDDREF 1701 1867 VDDREF pch l=0.04u w=0.8u
m17173 VDDREF 1702 1871 VDDREF pch l=0.04u w=0.8u
m17174 VDDREF 1906 29167 VDDREF pch l=0.04u w=0.12u
m17175 1880 1834 VDDREF VDDREF pch l=0.04u w=0.8u
m17176 1882 1835 VDDREF VDDREF pch l=0.04u w=0.8u
m17177 1884 1836 VDDREF VDDREF pch l=0.04u w=0.8u
m17178 1885 1837 VDDREF VDDREF pch l=0.04u w=0.8u
m17179 1886 1838 VDDREF VDDREF pch l=0.04u w=0.8u
m17180 1888 1839 VDDREF VDDREF pch l=0.04u w=0.8u
m17181 1889 1840 VDDREF VDDREF pch l=0.04u w=0.8u
m17182 1890 1841 VDDREF VDDREF pch l=0.04u w=0.8u
m17183 1892 1842 VDDREF VDDREF pch l=0.04u w=0.8u
m17184 1893 1843 VDDREF VDDREF pch l=0.04u w=0.8u
m17185 VDDREF FBDIV[5] 1875 VDDREF pch l=0.04u w=0.8u
m17186 1894 1934 VDDREF VDDREF pch l=0.04u w=0.8u
m17187 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m17188 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m17189 VDDREF 1983 1821 VDDREF pch l=0.04u w=0.8u
m17190 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m17191 VDDREF 1909 29173 VDDREF pch l=0.04u w=0.12u
m17192 VDDREF 1910 29174 VDDREF pch l=0.04u w=0.12u
m17193 1878 11 VDDREF VDDREF pch l=0.04u w=0.8u
m17194 1899 1917 29176 VDDREF pch l=0.04u w=0.12u
m17195 1895 1799 1863 VDDREF pch l=0.04u w=0.8u
m17196 1896 1800 1864 VDDREF pch l=0.04u w=0.8u
m17197 1897 1801 1865 VDDREF pch l=0.04u w=0.8u
m17198 1898 1802 1866 VDDREF pch l=0.04u w=0.8u
m17199 1906 1854 VDDREF VDDREF pch l=0.04u w=0.8u
m17200 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m17201 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m17202 1900 1807 1868 VDDREF pch l=0.04u w=0.8u
m17203 1901 1808 1869 VDDREF pch l=0.04u w=0.8u
m17204 1902 1809 1870 VDDREF pch l=0.04u w=0.8u
m17205 1879 979 VDDREF VDDREF pch l=0.04u w=0.8u
m17206 VDDREF 1720 1880 VDDREF pch l=0.04u w=0.8u
m17207 1881 1660 VDDREF VDDREF pch l=0.04u w=0.8u
m17208 VDDREF 1722 1882 VDDREF pch l=0.04u w=0.8u
m17209 1903 1810 1872 VDDREF pch l=0.04u w=0.8u
m17210 1904 1811 1873 VDDREF pch l=0.04u w=0.8u
m17211 1905 1812 1874 VDDREF pch l=0.04u w=0.8u
m17212 1883 1657 VDDREF VDDREF pch l=0.04u w=0.8u
m17213 VDDREF 1727 1884 VDDREF pch l=0.04u w=0.8u
m17214 VDDREF 1728 1885 VDDREF pch l=0.04u w=0.8u
m17215 VDDREF 1729 1886 VDDREF pch l=0.04u w=0.8u
m17216 1887 1577 VDDREF VDDREF pch l=0.04u w=0.8u
m17217 VDDREF 1731 1888 VDDREF pch l=0.04u w=0.8u
m17218 VDDREF 1732 1889 VDDREF pch l=0.04u w=0.8u
m17219 VDDREF 1733 1890 VDDREF pch l=0.04u w=0.8u
m17220 1891 1579 VDDREF VDDREF pch l=0.04u w=0.8u
m17221 VDDREF 1735 1892 VDDREF pch l=0.04u w=0.8u
m17222 VDDREF 1736 1893 VDDREF pch l=0.04u w=0.8u
m17223 1908 94 VDDREF VDDREF pch l=0.04u w=0.8u
m17224 1821 1983 VDDREF VDDREF pch l=0.04u w=0.8u
m17225 1909 1861 VDDREF VDDREF pch l=0.04u w=0.8u
m17226 1910 1862 VDDREF VDDREF pch l=0.04u w=0.8u
m17227 VDDREF 1976 1878 VDDREF pch l=0.04u w=0.8u
m17228 1911 3012 1899 VDDREF pch l=0.04u w=0.8u
m17229 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m17230 29188 4328 1895 VDDREF pch l=0.04u w=0.12u
m17231 29189 4328 1896 VDDREF pch l=0.04u w=0.12u
m17232 29190 4328 1897 VDDREF pch l=0.04u w=0.12u
m17233 29191 4328 1898 VDDREF pch l=0.04u w=0.12u
m17234 1912 1755 VDDREF VDDREF pch l=0.04u w=0.8u
m17235 29192 4328 1900 VDDREF pch l=0.04u w=0.12u
m17236 29193 4328 1901 VDDREF pch l=0.04u w=0.12u
m17237 29194 4328 1902 VDDREF pch l=0.04u w=0.12u
m17238 VDDREF 1657 1879 VDDREF pch l=0.04u w=0.8u
m17239 1913 1756 VDDREF VDDREF pch l=0.04u w=0.8u
m17240 VDDREF 139 1881 VDDREF pch l=0.04u w=0.8u
m17241 29195 4328 1903 VDDREF pch l=0.04u w=0.12u
m17242 29196 4328 1904 VDDREF pch l=0.04u w=0.12u
m17243 29197 4328 1905 VDDREF pch l=0.04u w=0.12u
m17244 VDDREF FRAC[19] 1883 VDDREF pch l=0.04u w=0.8u
m17245 VDDREF 1446 1887 VDDREF pch l=0.04u w=0.8u
m17246 VDDREF FRAC[19] 1891 VDDREF pch l=0.04u w=0.8u
m17247 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m17248 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m17249 1914 1850 VDDREF VDDREF pch l=0.04u w=0.8u
m17250 VDDREF 1934 1907 VDDREF pch l=0.04u w=0.8u
m17251 1915 377 VDDREF VDDREF pch l=0.04u w=0.8u
m17252 VDDREF 1936 1821 VDDREF pch l=0.04u w=0.8u
m17253 VDDREF 1937 VDDREF VDDREF pch l=0.26u w=1u
m17254 VDDREF 1941 29188 VDDREF pch l=0.04u w=0.12u
m17255 VDDREF 1505 29189 VDDREF pch l=0.04u w=0.12u
m17256 VDDREF 1942 29190 VDDREF pch l=0.04u w=0.12u
m17257 VDDREF 1508 29191 VDDREF pch l=0.04u w=0.12u
m17258 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m17259 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m17260 VDDREF 688 29192 VDDREF pch l=0.04u w=0.12u
m17261 VDDREF 1789 29193 VDDREF pch l=0.04u w=0.12u
m17262 VDDREF 731 29194 VDDREF pch l=0.04u w=0.12u
m17263 VDDREF 1943 29195 VDDREF pch l=0.04u w=0.12u
m17264 VDDREF 1791 29196 VDDREF pch l=0.04u w=0.12u
m17265 VDDREF 735 29197 VDDREF pch l=0.04u w=0.12u
m17266 1920 1774 VDDREF VDDREF pch l=0.04u w=0.8u
m17267 1922 1776 VDDREF VDDREF pch l=0.04u w=0.8u
m17268 1924 1778 VDDREF VDDREF pch l=0.04u w=0.8u
m17269 1925 1780 VDDREF VDDREF pch l=0.04u w=0.8u
m17270 1926 1781 VDDREF VDDREF pch l=0.04u w=0.8u
m17271 1928 1783 VDDREF VDDREF pch l=0.04u w=0.8u
m17272 1929 1784 VDDREF VDDREF pch l=0.04u w=0.8u
m17273 1930 1785 VDDREF VDDREF pch l=0.04u w=0.8u
m17274 1932 1787 VDDREF VDDREF pch l=0.04u w=0.8u
m17275 1933 1788 VDDREF VDDREF pch l=0.04u w=0.8u
m17276 VDDREF 1906 1914 VDDREF pch l=0.04u w=0.8u
m17277 1935 398 VDDREF VDDREF pch l=0.04u w=0.8u
m17278 1938 1938 VDDREF VDDREF pch l=0.04u w=1u
m17279 VDDREF 1952 VDDREF VDDREF pch l=0.26u w=1u
m17280 1939 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17281 1940 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17282 1941 1895 VDDREF VDDREF pch l=0.04u w=0.8u
m17283 1505 1896 VDDREF VDDREF pch l=0.04u w=0.8u
m17284 1942 1897 VDDREF VDDREF pch l=0.04u w=0.8u
m17285 1508 1898 VDDREF VDDREF pch l=0.04u w=0.8u
m17286 1916 303 VDDREF VDDREF pch l=0.04u w=0.8u
m17287 VDDREF 3012 1917 VDDREF pch l=0.04u w=0.8u
m17288 688 1900 VDDREF VDDREF pch l=0.04u w=0.8u
m17289 1789 1901 VDDREF VDDREF pch l=0.04u w=0.8u
m17290 VDDREF 1953 VDDREF VDDREF pch l=0.26u w=1u
m17291 731 1902 VDDREF VDDREF pch l=0.04u w=0.8u
m17292 1943 1903 VDDREF VDDREF pch l=0.04u w=0.8u
m17293 1791 1904 VDDREF VDDREF pch l=0.04u w=0.8u
m17294 VDDREF 1955 VDDREF VDDREF pch l=0.26u w=1u
m17295 735 1905 VDDREF VDDREF pch l=0.04u w=0.8u
m17296 1918 1581 1755 VDDREF pch l=0.04u w=0.8u
m17297 1819 1957 1919 VDDREF pch l=0.04u w=0.8u
m17298 458 1585 1756 VDDREF pch l=0.04u w=0.8u
m17299 1944 1958 1921 VDDREF pch l=0.04u w=0.8u
m17300 1946 1959 1923 VDDREF pch l=0.04u w=0.8u
m17301 1443 1960 1927 VDDREF pch l=0.04u w=0.8u
m17302 1445 1961 1931 VDDREF pch l=0.04u w=0.8u
m17303 1934 1982 VDDREF VDDREF pch l=0.04u w=0.8u
m17304 1948 377 VDDREF VDDREF pch l=0.04u w=0.8u
m17305 1936 2079 VDDREF VDDREF pch l=0.04u w=0.8u
m17306 1951 1951 VDDREF VDDREF pch l=0.04u w=1u
m17307 VDDREF 149 1916 VDDREF pch l=0.04u w=0.8u
m17308 VDDREF 1969 VDDREF VDDREF pch l=0.26u w=1u
m17309 VDDREF 1970 VDDREF VDDREF pch l=0.26u w=1u
m17310 1954 1954 VDDREF VDDREF pch l=0.04u w=1u
m17311 1956 1956 VDDREF VDDREF pch l=0.04u w=1u
m17312 1581 1755 1918 VDDREF pch l=0.04u w=0.8u
m17313 1957 1919 1819 VDDREF pch l=0.04u w=0.8u
m17314 1585 1756 458 VDDREF pch l=0.04u w=0.8u
m17315 1958 1921 1944 VDDREF pch l=0.04u w=0.8u
m17316 1959 1923 1946 VDDREF pch l=0.04u w=0.8u
m17317 1960 1927 1443 VDDREF pch l=0.04u w=0.8u
m17318 1961 1931 1445 VDDREF pch l=0.04u w=0.8u
m17319 1820 1594 1774 VDDREF pch l=0.04u w=0.8u
m17320 1945 1595 1776 VDDREF pch l=0.04u w=0.8u
m17321 1790 1596 1778 VDDREF pch l=0.04u w=0.8u
m17322 1770 1597 1780 VDDREF pch l=0.04u w=0.8u
m17323 1947 1598 1781 VDDREF pch l=0.04u w=0.8u
m17324 1626 1599 1783 VDDREF pch l=0.04u w=0.8u
m17325 1805 1600 1784 VDDREF pch l=0.04u w=0.8u
m17326 1793 1601 1785 VDDREF pch l=0.04u w=0.8u
m17327 1628 1602 1787 VDDREF pch l=0.04u w=0.8u
m17328 1806 1603 1788 VDDREF pch l=0.04u w=0.8u
m17329 1962 1914 VDDREF VDDREF pch l=0.04u w=0.8u
m17330 VDDREF 2648 1934 VDDREF pch l=0.04u w=0.8u
m17331 VDDREF REFDIV[3] 1948 VDDREF pch l=0.04u w=0.8u
m17332 VDDREF 2023 1936 VDDREF pch l=0.04u w=0.8u
m17333 1963 593 VDDREF VDDREF pch l=0.04u w=0.8u
m17334 VDDREF 1949 1950 VDDREF pch l=0.04u w=1u
m17335 1968 1968 VDDREF VDDREF pch l=0.04u w=1u
m17336 1971 1971 VDDREF VDDREF pch l=0.04u w=1u
m17337 1964 4328 1909 VDDREF pch l=0.04u w=0.8u
m17338 1965 4328 1910 VDDREF pch l=0.04u w=0.8u
m17339 1972 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17340 1973 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17341 1974 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17342 1975 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17343 1911 1593 VDDREF VDDREF pch l=0.04u w=0.8u
m17344 1594 1774 1820 VDDREF pch l=0.04u w=0.8u
m17345 1595 1776 1945 VDDREF pch l=0.04u w=0.8u
m17346 1596 1778 1790 VDDREF pch l=0.04u w=0.8u
m17347 1597 1780 1770 VDDREF pch l=0.04u w=0.8u
m17348 1598 1781 1947 VDDREF pch l=0.04u w=0.8u
m17349 1599 1783 1626 VDDREF pch l=0.04u w=0.8u
m17350 1600 1784 1805 VDDREF pch l=0.04u w=0.8u
m17351 1601 1785 1793 VDDREF pch l=0.04u w=0.8u
m17352 1602 1787 1628 VDDREF pch l=0.04u w=0.8u
m17353 1603 1788 1806 VDDREF pch l=0.04u w=0.8u
m17354 VDDREF 1875 1962 VDDREF pch l=0.04u w=0.8u
m17355 VDDREF 1967 1966 VDDREF pch l=0.04u w=1u
m17356 29238 1939 1964 VDDREF pch l=0.04u w=0.12u
m17357 29239 1940 1965 VDDREF pch l=0.04u w=0.12u
m17358 VDDREF 149 1976 VDDREF pch l=0.04u w=0.8u
m17359 VDDREF 1740 1911 VDDREF pch l=0.04u w=0.8u
m17360 1990 110 VDDREF VDDREF pch l=0.04u w=0.8u
m17361 VDDREF 1957 1977 VDDREF pch l=0.04u w=0.8u
m17362 1991 2022 VDDREF VDDREF pch l=0.04u w=0.8u
m17363 VDDREF 1958 1978 VDDREF pch l=0.04u w=0.8u
m17364 VDDREF 1959 1979 VDDREF pch l=0.04u w=0.8u
m17365 VDDREF 1960 1980 VDDREF pch l=0.04u w=0.8u
m17366 VDDREF 1961 1981 VDDREF pch l=0.04u w=0.8u
m17367 VDDREF 2021 1982 VDDREF pch l=0.04u w=0.8u
m17368 1997 1915 VDDREF VDDREF pch l=0.04u w=0.8u
m17369 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17370 1983 REFDIV[4] VDDREF VDDREF pch l=0.04u w=0.8u
m17371 1998 294 VDDREF VDDREF pch l=0.04u w=0.8u
m17372 VDDREF 2017 29238 VDDREF pch l=0.04u w=0.12u
m17373 VDDREF 2018 29239 VDDREF pch l=0.04u w=0.12u
m17374 VDDREF 1985 1984 VDDREF pch l=0.04u w=1u
m17375 VDDREF 1986 1987 VDDREF pch l=0.04u w=1u
m17376 1999 4328 1988 VDDREF pch l=0.04u w=0.8u
m17377 2000 4328 1947 VDDREF pch l=0.04u w=0.8u
m17378 2001 4328 1989 VDDREF pch l=0.04u w=0.8u
m17379 2002 4328 1793 VDDREF pch l=0.04u w=0.8u
m17380 VDDREF 592 1990 VDDREF pch l=0.04u w=0.8u
m17381 VDDREF 735 1991 VDDREF pch l=0.04u w=0.8u
m17382 VDDREF 1992 1993 VDDREF pch l=0.04u w=1u
m17383 2003 2073 VDDREF VDDREF pch l=0.04u w=0.8u
m17384 2004 2086 VDDREF VDDREF pch l=0.04u w=0.8u
m17385 2005 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m17386 2006 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m17387 VDDREF 1994 1995 VDDREF pch l=0.04u w=1u
m17388 2007 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m17389 2008 FRAC[6] VDDREF VDDREF pch l=0.04u w=0.8u
m17390 VDDREF 2053 1996 VDDREF pch l=0.04u w=0.8u
m17391 2009 2074 VDDREF VDDREF pch l=0.04u w=0.8u
m17392 2010 2088 VDDREF VDDREF pch l=0.04u w=0.8u
m17393 2011 1989 VDDREF VDDREF pch l=0.04u w=0.8u
m17394 2012 1996 VDDREF VDDREF pch l=0.04u w=0.8u
m17395 2013 2089 VDDREF VDDREF pch l=0.04u w=0.8u
m17396 2014 FRAC[6] VDDREF VDDREF pch l=0.04u w=0.8u
m17397 2015 1996 VDDREF VDDREF pch l=0.04u w=0.8u
m17398 29249 1907 VDDREF VDDREF pch l=0.04u w=0.24u
m17399 VDDREF 1860 1997 VDDREF pch l=0.04u w=0.8u
m17400 VDDREF 377 1983 VDDREF pch l=0.04u w=0.8u
m17401 2016 2016 VDDREF VDDREF pch l=0.04u w=1u
m17402 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17403 2017 1964 VDDREF VDDREF pch l=0.04u w=0.8u
m17404 2018 1965 VDDREF VDDREF pch l=0.04u w=0.8u
m17405 29255 1972 1999 VDDREF pch l=0.04u w=0.12u
m17406 29256 1973 2000 VDDREF pch l=0.04u w=0.12u
m17407 29257 1974 2001 VDDREF pch l=0.04u w=0.12u
m17408 29258 1975 2002 VDDREF pch l=0.04u w=0.12u
m17409 2019 3012 VDDREF VDDREF pch l=0.04u w=0.8u
m17410 2020 303 VDDREF VDDREF pch l=0.04u w=0.8u
m17411 1638 2158 VDDREF VDDREF pch l=0.04u w=0.8u
m17412 VDDREF 2071 2003 VDDREF pch l=0.04u w=0.8u
m17413 1640 2160 VDDREF VDDREF pch l=0.04u w=0.8u
m17414 VDDREF 2072 2004 VDDREF pch l=0.04u w=0.8u
m17415 VDDREF 2223 2005 VDDREF pch l=0.04u w=0.8u
m17416 VDDREF 2224 2006 VDDREF pch l=0.04u w=0.8u
m17417 VDDREF 596 2007 VDDREF pch l=0.04u w=0.8u
m17418 1642 2162 VDDREF VDDREF pch l=0.04u w=0.8u
m17419 VDDREF 2073 2008 VDDREF pch l=0.04u w=0.8u
m17420 VDDREF 131 2009 VDDREF pch l=0.04u w=0.8u
m17421 VDDREF 2074 2010 VDDREF pch l=0.04u w=0.8u
m17422 1646 2166 VDDREF VDDREF pch l=0.04u w=0.8u
m17423 VDDREF 2075 2011 VDDREF pch l=0.04u w=0.8u
m17424 VDDREF 2076 2012 VDDREF pch l=0.04u w=0.8u
m17425 VDDREF 2077 2013 VDDREF pch l=0.04u w=0.8u
m17426 1650 2170 VDDREF VDDREF pch l=0.04u w=0.8u
m17427 VDDREF 2078 2014 VDDREF pch l=0.04u w=0.8u
m17428 VDDREF FBDIV[6] 2015 VDDREF pch l=0.04u w=0.8u
m17429 2021 2188 29249 VDDREF pch l=0.04u w=0.24u
m17430 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17431 2024 129 VDDREF VDDREF pch l=0.04u w=0.8u
m17432 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17433 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17434 VDDREF 2034 29255 VDDREF pch l=0.04u w=0.12u
m17435 VDDREF 2035 29256 VDDREF pch l=0.04u w=0.12u
m17436 VDDREF 2036 29257 VDDREF pch l=0.04u w=0.12u
m17437 VDDREF 2037 29258 VDDREF pch l=0.04u w=0.12u
m17438 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17439 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17440 2027 592 VDDREF VDDREF pch l=0.04u w=0.8u
m17441 VDDREF 2055 1638 VDDREF pch l=0.04u w=0.8u
m17442 2028 735 VDDREF VDDREF pch l=0.04u w=0.8u
m17443 VDDREF 2057 1640 VDDREF pch l=0.04u w=0.8u
m17444 VDDREF 2059 1642 VDDREF pch l=0.04u w=0.8u
m17445 VDDREF 2064 1646 VDDREF pch l=0.04u w=0.8u
m17446 VDDREF 2068 1650 VDDREF pch l=0.04u w=0.8u
m17447 2029 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17448 2030 2151 2021 VDDREF pch l=0.04u w=0.8u
m17449 VDDREF 3454 2022 VDDREF pch l=0.04u w=0.8u
m17450 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17451 2031 1997 VDDREF VDDREF pch l=0.04u w=0.8u
m17452 VDDREF 377 2023 VDDREF pch l=0.04u w=0.8u
m17453 2032 1939 2017 VDDREF pch l=0.04u w=0.8u
m17454 2033 1940 2018 VDDREF pch l=0.04u w=0.8u
m17455 2034 1999 VDDREF VDDREF pch l=0.04u w=0.8u
m17456 2035 2000 VDDREF VDDREF pch l=0.04u w=0.8u
m17457 2036 2001 VDDREF VDDREF pch l=0.04u w=0.8u
m17458 2037 2002 VDDREF VDDREF pch l=0.04u w=0.8u
m17459 2025 2019 VDDREF VDDREF pch l=0.04u w=0.8u
m17460 2026 2020 VDDREF VDDREF pch l=0.04u w=0.8u
m17461 2040 2071 VDDREF VDDREF pch l=0.04u w=0.8u
m17462 2041 2072 VDDREF VDDREF pch l=0.04u w=0.8u
m17463 2042 2005 VDDREF VDDREF pch l=0.04u w=0.8u
m17464 2043 2006 VDDREF VDDREF pch l=0.04u w=0.8u
m17465 2044 2007 VDDREF VDDREF pch l=0.04u w=0.8u
m17466 2045 2073 VDDREF VDDREF pch l=0.04u w=0.8u
m17467 2046 131 VDDREF VDDREF pch l=0.04u w=0.8u
m17468 2047 2074 VDDREF VDDREF pch l=0.04u w=0.8u
m17469 2048 2075 VDDREF VDDREF pch l=0.04u w=0.8u
m17470 2049 2076 VDDREF VDDREF pch l=0.04u w=0.8u
m17471 2050 2077 VDDREF VDDREF pch l=0.04u w=0.8u
m17472 2051 2078 VDDREF VDDREF pch l=0.04u w=0.8u
m17473 2052 FBDIV[6] VDDREF VDDREF pch l=0.04u w=0.8u
m17474 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17475 VDDREF 1948 2031 VDDREF pch l=0.04u w=0.8u
m17476 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17477 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17478 2054 441 VDDREF VDDREF pch l=0.04u w=0.8u
m17479 29280 4328 2032 VDDREF pch l=0.04u w=0.12u
m17480 29281 4328 2033 VDDREF pch l=0.04u w=0.12u
m17481 VDDREF 2270 2025 VDDREF pch l=0.04u w=0.8u
m17482 VDDREF 2271 2026 VDDREF pch l=0.04u w=0.8u
m17483 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17484 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17485 2038 110 592 VDDREF pch l=0.04u w=0.8u
m17486 2055 1919 VDDREF VDDREF pch l=0.04u w=0.8u
m17487 2039 2022 735 VDDREF pch l=0.04u w=0.8u
m17488 2057 1921 VDDREF VDDREF pch l=0.04u w=0.8u
m17489 2059 1923 VDDREF VDDREF pch l=0.04u w=0.8u
m17490 2064 1927 VDDREF VDDREF pch l=0.04u w=0.8u
m17491 2068 1931 VDDREF VDDREF pch l=0.04u w=0.8u
m17492 2061 4328 2053 VDDREF pch l=0.04u w=0.8u
m17493 2030 2122 VDDREF VDDREF pch l=0.04u w=0.8u
m17494 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17495 2031 1948 VDDREF VDDREF pch l=0.04u w=0.8u
m17496 VDDREF 60 29280 VDDREF pch l=0.04u w=0.12u
m17497 VDDREF 2098 29281 VDDREF pch l=0.04u w=0.12u
m17498 2080 1972 2034 VDDREF pch l=0.04u w=0.8u
m17499 2081 1973 2035 VDDREF pch l=0.04u w=0.8u
m17500 2082 1974 2036 VDDREF pch l=0.04u w=0.8u
m17501 2083 1975 2037 VDDREF pch l=0.04u w=0.8u
m17502 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17503 110 592 2038 VDDREF pch l=0.04u w=0.8u
m17504 VDDREF 1957 2055 VDDREF pch l=0.04u w=0.8u
m17505 2022 735 2039 VDDREF pch l=0.04u w=0.8u
m17506 VDDREF 1958 2057 VDDREF pch l=0.04u w=0.8u
m17507 VDDREF 1959 2059 VDDREF pch l=0.04u w=0.8u
m17508 VDDREF 1960 2064 VDDREF pch l=0.04u w=0.8u
m17509 VDDREF 1961 2068 VDDREF pch l=0.04u w=0.8u
m17510 2090 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17511 2091 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17512 2092 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17513 2056 2073 2071 VDDREF pch l=0.04u w=0.8u
m17514 2058 2086 2072 VDDREF pch l=0.04u w=0.8u
m17515 2093 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17516 2094 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17517 2095 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17518 2060 FRAC[6] 2073 VDDREF pch l=0.04u w=0.8u
m17519 29292 2029 2061 VDDREF pch l=0.04u w=0.12u
m17520 2062 2074 131 VDDREF pch l=0.04u w=0.8u
m17521 2063 2088 2074 VDDREF pch l=0.04u w=0.8u
m17522 2065 1989 2075 VDDREF pch l=0.04u w=0.8u
m17523 2066 1996 2076 VDDREF pch l=0.04u w=0.8u
m17524 2067 2089 2077 VDDREF pch l=0.04u w=0.8u
m17525 2069 FRAC[6] 2078 VDDREF pch l=0.04u w=0.8u
m17526 2070 1996 FBDIV[6] VDDREF pch l=0.04u w=0.8u
m17527 VDDREF 2648 2030 VDDREF pch l=0.04u w=0.8u
m17528 VDDREF 1997 2031 VDDREF pch l=0.04u w=0.8u
m17529 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17530 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17531 2079 2104 1677 VDDREF pch l=0.04u w=0.8u
m17532 2097 735 VDDREF VDDREF pch l=0.04u w=0.8u
m17533 60 2032 VDDREF VDDREF pch l=0.04u w=0.8u
m17534 2098 2033 VDDREF VDDREF pch l=0.04u w=0.8u
m17535 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17536 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17537 29296 4328 2080 VDDREF pch l=0.04u w=0.12u
m17538 29297 4328 2081 VDDREF pch l=0.04u w=0.12u
m17539 29298 4328 2082 VDDREF pch l=0.04u w=0.12u
m17540 29299 4328 2083 VDDREF pch l=0.04u w=0.12u
m17541 VDDREF 4353 2084 VDDREF pch l=0.04u w=0.8u
m17542 VDDREF 11 2085 VDDREF pch l=0.04u w=0.8u
m17543 2073 2071 2056 VDDREF pch l=0.04u w=0.8u
m17544 2086 2072 2058 VDDREF pch l=0.04u w=0.8u
m17545 FRAC[6] 2073 2060 VDDREF pch l=0.04u w=0.8u
m17546 VDDREF 2111 29292 VDDREF pch l=0.04u w=0.12u
m17547 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17548 2074 131 2062 VDDREF pch l=0.04u w=0.8u
m17549 2088 2074 2063 VDDREF pch l=0.04u w=0.8u
m17550 1989 2075 2065 VDDREF pch l=0.04u w=0.8u
m17551 1996 2076 2066 VDDREF pch l=0.04u w=0.8u
m17552 2089 2077 2067 VDDREF pch l=0.04u w=0.8u
m17553 FRAC[6] 2078 2069 VDDREF pch l=0.04u w=0.8u
m17554 1996 FBDIV[6] 2070 VDDREF pch l=0.04u w=0.8u
m17555 29304 2030 VDDREF VDDREF pch l=0.04u w=0.12u
m17556 2104 1677 2079 VDDREF pch l=0.04u w=0.8u
m17557 VDDREF 2075 29296 VDDREF pch l=0.04u w=0.12u
m17558 VDDREF 1792 29297 VDDREF pch l=0.04u w=0.12u
m17559 VDDREF 2078 29298 VDDREF pch l=0.04u w=0.12u
m17560 VDDREF 1794 29299 VDDREF pch l=0.04u w=0.12u
m17561 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17562 2099 2038 VDDREF VDDREF pch l=0.04u w=0.8u
m17563 1957 688 1943 VDDREF pch l=0.04u w=0.8u
m17564 2100 2039 VDDREF VDDREF pch l=0.04u w=0.8u
m17565 1958 1946 139 VDDREF pch l=0.04u w=0.8u
m17566 1959 1943 FRAC[18] VDDREF pch l=0.04u w=0.8u
m17567 2111 2061 VDDREF VDDREF pch l=0.04u w=0.8u
m17568 1960 1576 1445 VDDREF pch l=0.04u w=0.8u
m17569 1961 1578 FRAC[18] VDDREF pch l=0.04u w=0.8u
m17570 2122 2151 29304 VDDREF pch l=0.04u w=0.12u
m17571 2105 4328 2102 VDDREF pch l=0.04u w=0.8u
m17572 2106 4328 2103 VDDREF pch l=0.04u w=0.8u
m17573 2107 4328 595 VDDREF pch l=0.04u w=0.8u
m17574 2108 4328 2042 VDDREF pch l=0.04u w=0.8u
m17575 2109 4328 2043 VDDREF pch l=0.04u w=0.8u
m17576 2110 4328 2044 VDDREF pch l=0.04u w=0.8u
m17577 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17578 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17579 2123 76 VDDREF VDDREF pch l=0.04u w=0.8u
m17580 VDDREF 2096 2104 VDDREF pch l=0.04u w=0.8u
m17581 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17582 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17583 139 1027 VDDREF VDDREF pch l=0.04u w=0.8u
m17584 2124 2131 VDDREF VDDREF pch l=0.04u w=0.8u
m17585 2125 1099 VDDREF VDDREF pch l=0.04u w=0.8u
m17586 2075 2080 VDDREF VDDREF pch l=0.04u w=0.8u
m17587 1792 2081 VDDREF VDDREF pch l=0.04u w=0.8u
m17588 2078 2082 VDDREF VDDREF pch l=0.04u w=0.8u
m17589 1794 2083 VDDREF VDDREF pch l=0.04u w=0.8u
m17590 2126 4353 2025 VDDREF pch l=0.04u w=0.8u
m17591 2127 11 2026 VDDREF pch l=0.04u w=0.8u
m17592 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17593 VDDREF 1867 2099 VDDREF pch l=0.04u w=0.8u
m17594 688 1943 1957 VDDREF pch l=0.04u w=0.8u
m17595 VDDREF 1871 2100 VDDREF pch l=0.04u w=0.8u
m17596 1946 139 1958 VDDREF pch l=0.04u w=0.8u
m17597 1943 FRAC[18] 1959 VDDREF pch l=0.04u w=0.8u
m17598 1576 1445 1960 VDDREF pch l=0.04u w=0.8u
m17599 1578 FRAC[18] 1961 VDDREF pch l=0.04u w=0.8u
m17600 1934 2188 2122 VDDREF pch l=0.04u w=0.8u
m17601 29318 2090 2105 VDDREF pch l=0.04u w=0.12u
m17602 29319 2091 2106 VDDREF pch l=0.04u w=0.12u
m17603 29320 2092 2107 VDDREF pch l=0.04u w=0.12u
m17604 2112 2056 VDDREF VDDREF pch l=0.04u w=0.8u
m17605 2113 2058 VDDREF VDDREF pch l=0.04u w=0.8u
m17606 29321 2093 2108 VDDREF pch l=0.04u w=0.12u
m17607 29322 2094 2109 VDDREF pch l=0.04u w=0.12u
m17608 29323 2095 2110 VDDREF pch l=0.04u w=0.12u
m17609 2114 2060 VDDREF VDDREF pch l=0.04u w=0.8u
m17610 2115 2062 VDDREF VDDREF pch l=0.04u w=0.8u
m17611 2116 2063 VDDREF VDDREF pch l=0.04u w=0.8u
m17612 2117 2065 VDDREF VDDREF pch l=0.04u w=0.8u
m17613 2118 2066 VDDREF VDDREF pch l=0.04u w=0.8u
m17614 2119 2067 VDDREF VDDREF pch l=0.04u w=0.8u
m17615 2120 2069 VDDREF VDDREF pch l=0.04u w=0.8u
m17616 2121 2070 VDDREF VDDREF pch l=0.04u w=0.8u
m17617 2128 155 VDDREF VDDREF pch l=0.04u w=0.8u
m17618 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17619 29325 2084 2126 VDDREF pch l=0.04u w=0.12u
m17620 29326 2085 2127 VDDREF pch l=0.04u w=0.12u
m17621 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17622 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17623 VDDREF 2144 29318 VDDREF pch l=0.04u w=0.12u
m17624 VDDREF 2145 29319 VDDREF pch l=0.04u w=0.12u
m17625 VDDREF 2146 29320 VDDREF pch l=0.04u w=0.12u
m17626 VDDREF 1880 2112 VDDREF pch l=0.04u w=0.8u
m17627 VDDREF 1882 2113 VDDREF pch l=0.04u w=0.8u
m17628 VDDREF 2148 29321 VDDREF pch l=0.04u w=0.12u
m17629 VDDREF 2149 29322 VDDREF pch l=0.04u w=0.12u
m17630 VDDREF 2150 29323 VDDREF pch l=0.04u w=0.12u
m17631 VDDREF 1884 2114 VDDREF pch l=0.04u w=0.8u
m17632 2132 2029 2111 VDDREF pch l=0.04u w=0.8u
m17633 VDDREF 1885 2115 VDDREF pch l=0.04u w=0.8u
m17634 VDDREF 1886 2116 VDDREF pch l=0.04u w=0.8u
m17635 VDDREF 1888 2117 VDDREF pch l=0.04u w=0.8u
m17636 VDDREF 1889 2118 VDDREF pch l=0.04u w=0.8u
m17637 VDDREF 1890 2119 VDDREF pch l=0.04u w=0.8u
m17638 VDDREF 1892 2120 VDDREF pch l=0.04u w=0.8u
m17639 VDDREF 1893 2121 VDDREF pch l=0.04u w=0.8u
m17640 2138 76 2031 VDDREF pch l=0.04u w=0.8u
m17641 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17642 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17643 VDDREF 683 2096 VDDREF pch l=0.04u w=0.8u
m17644 140 3338 VDDREF VDDREF pch l=0.04u w=0.8u
m17645 2129 60 2131 VDDREF pch l=0.04u w=0.8u
m17646 2130 2098 1099 VDDREF pch l=0.04u w=0.8u
m17647 2139 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17648 2140 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17649 2141 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17650 2142 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17651 VDDREF 2156 29325 VDDREF pch l=0.04u w=0.12u
m17652 VDDREF 2157 29326 VDDREF pch l=0.04u w=0.12u
m17653 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17654 2143 2099 VDDREF VDDREF pch l=0.04u w=0.8u
m17655 2144 2105 VDDREF VDDREF pch l=0.04u w=0.8u
m17656 2145 2106 VDDREF VDDREF pch l=0.04u w=0.8u
m17657 2146 2107 VDDREF VDDREF pch l=0.04u w=0.8u
m17658 VDDREF 688 2133 VDDREF pch l=0.04u w=0.8u
m17659 2147 2100 VDDREF VDDREF pch l=0.04u w=0.8u
m17660 VDDREF 1946 2134 VDDREF pch l=0.04u w=0.8u
m17661 2148 2108 VDDREF VDDREF pch l=0.04u w=0.8u
m17662 2149 2109 VDDREF VDDREF pch l=0.04u w=0.8u
m17663 2150 2110 VDDREF VDDREF pch l=0.04u w=0.8u
m17664 VDDREF 1943 2135 VDDREF pch l=0.04u w=0.8u
m17665 29337 4328 2132 VDDREF pch l=0.04u w=0.12u
m17666 VDDREF 1576 2136 VDDREF pch l=0.04u w=0.8u
m17667 VDDREF 1578 2137 VDDREF pch l=0.04u w=0.8u
m17668 2151 2188 VDDREF VDDREF pch l=0.04u w=0.8u
m17669 2152 155 VDDREF VDDREF pch l=0.04u w=0.8u
m17670 29338 2123 2138 VDDREF pch l=0.04u w=0.12u
m17671 2096 1240 VDDREF VDDREF pch l=0.04u w=0.8u
m17672 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17673 60 2131 2129 VDDREF pch l=0.04u w=0.8u
m17674 2098 1099 2130 VDDREF pch l=0.04u w=0.8u
m17675 2156 2716 VDDREF VDDREF pch l=0.04u w=0.8u
m17676 2157 2716 VDDREF VDDREF pch l=0.04u w=0.8u
m17677 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17678 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17679 VDDREF 1990 2143 VDDREF pch l=0.04u w=0.8u
m17680 VDDREF 1991 2147 VDDREF pch l=0.04u w=0.8u
m17681 VDDREF 2184 29337 VDDREF pch l=0.04u w=0.12u
m17682 2159 2112 VDDREF VDDREF pch l=0.04u w=0.8u
m17683 2161 2113 VDDREF VDDREF pch l=0.04u w=0.8u
m17684 2163 2114 VDDREF VDDREF pch l=0.04u w=0.8u
m17685 2164 2115 VDDREF VDDREF pch l=0.04u w=0.8u
m17686 2165 2116 VDDREF VDDREF pch l=0.04u w=0.8u
m17687 2167 2117 VDDREF VDDREF pch l=0.04u w=0.8u
m17688 2168 2118 VDDREF VDDREF pch l=0.04u w=0.8u
m17689 2169 2119 VDDREF VDDREF pch l=0.04u w=0.8u
m17690 2171 2120 VDDREF VDDREF pch l=0.04u w=0.8u
m17691 2172 2121 VDDREF VDDREF pch l=0.04u w=0.8u
m17692 VDDREF FBDIV[6] 2152 VDDREF pch l=0.04u w=0.8u
m17693 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17694 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17695 VDDREF 2185 29338 VDDREF pch l=0.04u w=0.12u
m17696 VDDREF 2194 2096 VDDREF pch l=0.04u w=0.8u
m17697 459 3610 VDDREF VDDREF pch l=0.04u w=0.8u
m17698 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17699 2174 4328 2153 VDDREF pch l=0.04u w=0.8u
m17700 2175 4328 2154 VDDREF pch l=0.04u w=0.8u
m17701 2176 4328 2155 VDDREF pch l=0.04u w=0.8u
m17702 2177 4328 2076 VDDREF pch l=0.04u w=0.8u
m17703 VDDREF 2126 2156 VDDREF pch l=0.04u w=0.8u
m17704 VDDREF 2127 2157 VDDREF pch l=0.04u w=0.8u
m17705 2184 2132 VDDREF VDDREF pch l=0.04u w=0.8u
m17706 2178 2090 2144 VDDREF pch l=0.04u w=0.8u
m17707 2179 2091 2145 VDDREF pch l=0.04u w=0.8u
m17708 2180 2092 2146 VDDREF pch l=0.04u w=0.8u
m17709 2158 688 VDDREF VDDREF pch l=0.04u w=0.8u
m17710 VDDREF 2003 2159 VDDREF pch l=0.04u w=0.8u
m17711 2160 1946 VDDREF VDDREF pch l=0.04u w=0.8u
m17712 VDDREF 2004 2161 VDDREF pch l=0.04u w=0.8u
m17713 2181 2093 2148 VDDREF pch l=0.04u w=0.8u
m17714 2182 2094 2149 VDDREF pch l=0.04u w=0.8u
m17715 2183 2095 2150 VDDREF pch l=0.04u w=0.8u
m17716 2162 1943 VDDREF VDDREF pch l=0.04u w=0.8u
m17717 VDDREF 2008 2163 VDDREF pch l=0.04u w=0.8u
m17718 VDDREF 2009 2164 VDDREF pch l=0.04u w=0.8u
m17719 VDDREF 2010 2165 VDDREF pch l=0.04u w=0.8u
m17720 2166 1576 VDDREF VDDREF pch l=0.04u w=0.8u
m17721 VDDREF 2011 2167 VDDREF pch l=0.04u w=0.8u
m17722 VDDREF 2012 2168 VDDREF pch l=0.04u w=0.8u
m17723 VDDREF 2013 2169 VDDREF pch l=0.04u w=0.8u
m17724 2170 1578 VDDREF VDDREF pch l=0.04u w=0.8u
m17725 VDDREF 2014 2171 VDDREF pch l=0.04u w=0.8u
m17726 VDDREF 2015 2172 VDDREF pch l=0.04u w=0.8u
m17727 VDDREF 2188 2173 VDDREF pch l=0.04u w=0.8u
m17728 2185 2138 VDDREF VDDREF pch l=0.04u w=0.8u
m17729 VDDREF 2190 VDDREF VDDREF pch l=0.26u w=1u
m17730 29385 2139 2174 VDDREF pch l=0.04u w=0.12u
m17731 29386 2140 2175 VDDREF pch l=0.04u w=0.12u
m17732 29387 2141 2176 VDDREF pch l=0.04u w=0.12u
m17733 29388 2142 2177 VDDREF pch l=0.04u w=0.12u
m17734 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17735 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17736 2186 2038 VDDREF VDDREF pch l=0.04u w=0.8u
m17737 29543 4328 2178 VDDREF pch l=0.04u w=0.12u
m17738 29544 4328 2179 VDDREF pch l=0.04u w=0.12u
m17739 29545 4328 2180 VDDREF pch l=0.04u w=0.12u
m17740 VDDREF 1943 2158 VDDREF pch l=0.04u w=0.8u
m17741 2187 2039 VDDREF VDDREF pch l=0.04u w=0.8u
m17742 VDDREF 139 2160 VDDREF pch l=0.04u w=0.8u
m17743 29546 4328 2181 VDDREF pch l=0.04u w=0.12u
m17744 29547 4328 2182 VDDREF pch l=0.04u w=0.12u
m17745 29548 4328 2183 VDDREF pch l=0.04u w=0.12u
m17746 VDDREF FRAC[18] 2162 VDDREF pch l=0.04u w=0.8u
m17747 VDDREF 1445 2166 VDDREF pch l=0.04u w=0.8u
m17748 VDDREF FRAC[18] 2170 VDDREF pch l=0.04u w=0.8u
m17749 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17750 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17751 2189 2128 VDDREF VDDREF pch l=0.04u w=0.8u
m17752 2191 2191 VDDREF VDDREF pch l=0.04u w=1u
m17753 2192 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17754 2193 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17755 2194 2228 VDDREF VDDREF pch l=0.04u w=0.8u
m17756 VDDREF 2217 VDDREF VDDREF pch l=0.26u w=1u
m17757 VDDREF 2218 29385 VDDREF pch l=0.04u w=0.12u
m17758 VDDREF 2219 29386 VDDREF pch l=0.04u w=0.12u
m17759 VDDREF 2220 29387 VDDREF pch l=0.04u w=0.12u
m17760 VDDREF 2221 29388 VDDREF pch l=0.04u w=0.12u
m17761 755 3760 VDDREF VDDREF pch l=0.04u w=0.8u
m17762 2195 2084 2156 VDDREF pch l=0.04u w=0.8u
m17763 2196 2085 2157 VDDREF pch l=0.04u w=0.8u
m17764 VDDREF 395 29543 VDDREF pch l=0.04u w=0.12u
m17765 VDDREF 2071 29544 VDDREF pch l=0.04u w=0.12u
m17766 VDDREF 437 29545 VDDREF pch l=0.04u w=0.12u
m17767 VDDREF 2222 29546 VDDREF pch l=0.04u w=0.12u
m17768 VDDREF 2073 29547 VDDREF pch l=0.04u w=0.12u
m17769 VDDREF 441 29548 VDDREF pch l=0.04u w=0.12u
m17770 2199 2056 VDDREF VDDREF pch l=0.04u w=0.8u
m17771 2201 2058 VDDREF VDDREF pch l=0.04u w=0.8u
m17772 2203 2060 VDDREF VDDREF pch l=0.04u w=0.8u
m17773 2204 2062 VDDREF VDDREF pch l=0.04u w=0.8u
m17774 2205 2063 VDDREF VDDREF pch l=0.04u w=0.8u
m17775 2207 2065 VDDREF VDDREF pch l=0.04u w=0.8u
m17776 2208 2066 VDDREF VDDREF pch l=0.04u w=0.8u
m17777 2209 2067 VDDREF VDDREF pch l=0.04u w=0.8u
m17778 2211 2069 VDDREF VDDREF pch l=0.04u w=0.8u
m17779 2212 2070 VDDREF VDDREF pch l=0.04u w=0.8u
m17780 2188 2244 VDDREF VDDREF pch l=0.04u w=0.8u
m17781 VDDREF 2184 2189 VDDREF pch l=0.04u w=0.8u
m17782 2213 2123 2185 VDDREF pch l=0.04u w=0.8u
m17783 VDDREF 2228 2194 VDDREF pch l=0.04u w=0.8u
m17784 2216 2216 VDDREF VDDREF pch l=0.04u w=1u
m17785 2218 2174 VDDREF VDDREF pch l=0.04u w=0.8u
m17786 2219 2175 VDDREF VDDREF pch l=0.04u w=0.8u
m17787 2220 2176 VDDREF VDDREF pch l=0.04u w=0.8u
m17788 2221 2177 VDDREF VDDREF pch l=0.04u w=0.8u
m17789 VDDREF 2232 VDDREF VDDREF pch l=0.26u w=1u
m17790 VDDREF 2233 VDDREF VDDREF pch l=0.26u w=1u
m17791 29704 4353 2195 VDDREF pch l=0.04u w=0.24u
m17792 29705 11 2196 VDDREF pch l=0.04u w=0.24u
m17793 395 2178 VDDREF VDDREF pch l=0.04u w=0.8u
m17794 2071 2179 VDDREF VDDREF pch l=0.04u w=0.8u
m17795 VDDREF 2235 VDDREF VDDREF pch l=0.26u w=1u
m17796 437 2180 VDDREF VDDREF pch l=0.04u w=0.8u
m17797 2222 2181 VDDREF VDDREF pch l=0.04u w=0.8u
m17798 2073 2182 VDDREF VDDREF pch l=0.04u w=0.8u
m17799 VDDREF 2237 VDDREF VDDREF pch l=0.26u w=1u
m17800 441 2183 VDDREF VDDREF pch l=0.04u w=0.8u
m17801 2197 1867 2038 VDDREF pch l=0.04u w=0.8u
m17802 2102 2239 2198 VDDREF pch l=0.04u w=0.8u
m17803 754 1871 2039 VDDREF pch l=0.04u w=0.8u
m17804 2223 2240 2200 VDDREF pch l=0.04u w=0.8u
m17805 2225 2241 2202 VDDREF pch l=0.04u w=0.8u
m17806 1814 2242 2206 VDDREF pch l=0.04u w=0.8u
m17807 1815 2243 2210 VDDREF pch l=0.04u w=0.8u
m17808 VDDREF 2648 2188 VDDREF pch l=0.04u w=0.8u
m17809 29715 76 2213 VDDREF pch l=0.04u w=0.12u
m17810 VDDREF 2214 2215 VDDREF pch l=0.04u w=1u
m17811 2226 4328 2129 VDDREF pch l=0.04u w=0.8u
m17812 2227 4328 2130 VDDREF pch l=0.04u w=0.8u
m17813 2231 2231 VDDREF VDDREF pch l=0.04u w=1u
m17814 2234 2234 VDDREF VDDREF pch l=0.04u w=1u
m17815 VDDREF 2300 29704 VDDREF pch l=0.04u w=0.24u
m17816 VDDREF 2301 29705 VDDREF pch l=0.04u w=0.24u
m17817 1042 3479 VDDREF VDDREF pch l=0.04u w=0.8u
m17818 2236 2236 VDDREF VDDREF pch l=0.04u w=1u
m17819 2238 2238 VDDREF VDDREF pch l=0.04u w=1u
m17820 1867 2038 2197 VDDREF pch l=0.04u w=0.8u
m17821 2239 2198 2102 VDDREF pch l=0.04u w=0.8u
m17822 1871 2039 754 VDDREF pch l=0.04u w=0.8u
m17823 2240 2200 2223 VDDREF pch l=0.04u w=0.8u
m17824 2241 2202 2225 VDDREF pch l=0.04u w=0.8u
m17825 2242 2206 1814 VDDREF pch l=0.04u w=0.8u
m17826 2243 2210 1815 VDDREF pch l=0.04u w=0.8u
m17827 2103 1880 2056 VDDREF pch l=0.04u w=0.8u
m17828 2224 1882 2058 VDDREF pch l=0.04u w=0.8u
m17829 2072 1884 2060 VDDREF pch l=0.04u w=0.8u
m17830 2053 1885 2062 VDDREF pch l=0.04u w=0.8u
m17831 2154 1886 2063 VDDREF pch l=0.04u w=0.8u
m17832 1988 1888 2065 VDDREF pch l=0.04u w=0.8u
m17833 2088 1889 2066 VDDREF pch l=0.04u w=0.8u
m17834 2076 1890 2067 VDDREF pch l=0.04u w=0.8u
m17835 1989 1892 2069 VDDREF pch l=0.04u w=0.8u
m17836 2089 1893 2070 VDDREF pch l=0.04u w=0.8u
m17837 2245 2189 VDDREF VDDREF pch l=0.04u w=0.8u
m17838 VDDREF 1876 29715 VDDREF pch l=0.04u w=0.12u
m17839 29730 2192 2226 VDDREF pch l=0.04u w=0.12u
m17840 29731 2193 2227 VDDREF pch l=0.04u w=0.12u
m17841 2228 1742 VDDREF VDDREF pch l=0.04u w=0.8u
m17842 VDDREF 2230 2229 VDDREF pch l=0.04u w=1u
m17843 2246 2139 2218 VDDREF pch l=0.04u w=0.8u
m17844 2247 2140 2219 VDDREF pch l=0.04u w=0.8u
m17845 2248 2141 2220 VDDREF pch l=0.04u w=0.8u
m17846 2249 2142 2221 VDDREF pch l=0.04u w=0.8u
m17847 2250 2195 VDDREF VDDREF pch l=0.04u w=0.8u
m17848 2251 2196 VDDREF VDDREF pch l=0.04u w=0.8u
m17849 1880 2056 2103 VDDREF pch l=0.04u w=0.8u
m17850 1882 2058 2224 VDDREF pch l=0.04u w=0.8u
m17851 1884 2060 2072 VDDREF pch l=0.04u w=0.8u
m17852 1885 2062 2053 VDDREF pch l=0.04u w=0.8u
m17853 1886 2063 2154 VDDREF pch l=0.04u w=0.8u
m17854 1888 2065 1988 VDDREF pch l=0.04u w=0.8u
m17855 1889 2066 2088 VDDREF pch l=0.04u w=0.8u
m17856 1890 2067 2076 VDDREF pch l=0.04u w=0.8u
m17857 1892 2069 1989 VDDREF pch l=0.04u w=0.8u
m17858 1893 2070 2089 VDDREF pch l=0.04u w=0.8u
m17859 VDDREF 2285 2244 VDDREF pch l=0.04u w=0.8u
m17860 VDDREF 2152 2245 VDDREF pch l=0.04u w=0.8u
m17861 1876 2213 VDDREF VDDREF pch l=0.04u w=0.8u
m17862 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m17863 VDDREF 2268 29730 VDDREF pch l=0.04u w=0.12u
m17864 VDDREF 2269 29731 VDDREF pch l=0.04u w=0.12u
m17865 VDDREF 2286 2228 VDDREF pch l=0.04u w=0.8u
m17866 29773 4328 2246 VDDREF pch l=0.04u w=0.12u
m17867 29774 4328 2247 VDDREF pch l=0.04u w=0.12u
m17868 29775 4328 2248 VDDREF pch l=0.04u w=0.12u
m17869 29776 4328 2249 VDDREF pch l=0.04u w=0.12u
m17870 VDDREF 2253 2252 VDDREF pch l=0.04u w=1u
m17871 VDDREF 2254 2255 VDDREF pch l=0.04u w=1u
m17872 1514 3204 VDDREF VDDREF pch l=0.04u w=0.8u
m17873 2261 110 VDDREF VDDREF pch l=0.04u w=0.8u
m17874 VDDREF 2239 2256 VDDREF pch l=0.04u w=0.8u
m17875 2262 2290 VDDREF VDDREF pch l=0.04u w=0.8u
m17876 VDDREF 2240 2257 VDDREF pch l=0.04u w=0.8u
m17877 VDDREF 2241 2258 VDDREF pch l=0.04u w=0.8u
m17878 VDDREF 2242 2259 VDDREF pch l=0.04u w=0.8u
m17879 VDDREF 2243 2260 VDDREF pch l=0.04u w=0.8u
m17880 29932 2173 VDDREF VDDREF pch l=0.04u w=0.24u
m17881 2268 2226 VDDREF VDDREF pch l=0.04u w=0.8u
m17882 2269 2227 VDDREF VDDREF pch l=0.04u w=0.8u
m17883 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m17884 VDDREF 2287 29773 VDDREF pch l=0.04u w=0.12u
m17885 VDDREF 2074 29774 VDDREF pch l=0.04u w=0.12u
m17886 VDDREF 2288 29775 VDDREF pch l=0.04u w=0.12u
m17887 VDDREF 2077 29776 VDDREF pch l=0.04u w=0.12u
m17888 2270 2716 VDDREF VDDREF pch l=0.04u w=0.8u
m17889 2271 2716 VDDREF VDDREF pch l=0.04u w=0.8u
m17890 VDDREF 292 2261 VDDREF pch l=0.04u w=0.8u
m17891 VDDREF 1027 2262 VDDREF pch l=0.04u w=0.8u
m17892 2285 2454 29932 VDDREF pch l=0.04u w=0.24u
m17893 VDDREF 2263 2264 VDDREF pch l=0.04u w=1u
m17894 2272 2344 VDDREF VDDREF pch l=0.04u w=0.8u
m17895 2273 2357 VDDREF VDDREF pch l=0.04u w=0.8u
m17896 2274 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m17897 2275 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m17898 VDDREF 2265 2266 VDDREF pch l=0.04u w=1u
m17899 2276 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m17900 2277 FRAC[7] VDDREF VDDREF pch l=0.04u w=0.8u
m17901 VDDREF 2321 2267 VDDREF pch l=0.04u w=0.8u
m17902 2278 2345 VDDREF VDDREF pch l=0.04u w=0.8u
m17903 2279 2359 VDDREF VDDREF pch l=0.04u w=0.8u
m17904 2280 2324 VDDREF VDDREF pch l=0.04u w=0.8u
m17905 2281 2267 VDDREF VDDREF pch l=0.04u w=0.8u
m17906 2282 2360 VDDREF VDDREF pch l=0.04u w=0.8u
m17907 2283 FRAC[7] VDDREF VDDREF pch l=0.04u w=0.8u
m17908 2284 2267 VDDREF VDDREF pch l=0.04u w=0.8u
m17909 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m17910 2286 1876 VDDREF VDDREF pch l=0.04u w=0.8u
m17911 VDDREF 2400 VDDREF VDDREF pch l=0.26u w=1u
m17912 VDDREF 2401 VDDREF VDDREF pch l=0.26u w=1u
m17913 2287 2246 VDDREF VDDREF pch l=0.04u w=0.8u
m17914 2074 2247 VDDREF VDDREF pch l=0.04u w=0.8u
m17915 2288 2248 VDDREF VDDREF pch l=0.04u w=0.8u
m17916 2077 2249 VDDREF VDDREF pch l=0.04u w=0.8u
m17917 VDDREF 2250 2270 VDDREF pch l=0.04u w=0.8u
m17918 VDDREF 2251 2271 VDDREF pch l=0.04u w=0.8u
m17919 1803 2925 VDDREF VDDREF pch l=0.04u w=0.8u
m17920 2289 2403 2285 VDDREF pch l=0.04u w=0.8u
m17921 1919 2428 VDDREF VDDREF pch l=0.04u w=0.8u
m17922 VDDREF 2342 2272 VDDREF pch l=0.04u w=0.8u
m17923 1921 2430 VDDREF VDDREF pch l=0.04u w=0.8u
m17924 VDDREF 2343 2273 VDDREF pch l=0.04u w=0.8u
m17925 VDDREF 2488 2274 VDDREF pch l=0.04u w=0.8u
m17926 VDDREF 2489 2275 VDDREF pch l=0.04u w=0.8u
m17927 VDDREF 297 2276 VDDREF pch l=0.04u w=0.8u
m17928 1923 2432 VDDREF VDDREF pch l=0.04u w=0.8u
m17929 VDDREF 2344 2277 VDDREF pch l=0.04u w=0.8u
m17930 VDDREF 131 2278 VDDREF pch l=0.04u w=0.8u
m17931 VDDREF 2345 2279 VDDREF pch l=0.04u w=0.8u
m17932 1927 2436 VDDREF VDDREF pch l=0.04u w=0.8u
m17933 VDDREF 2346 2280 VDDREF pch l=0.04u w=0.8u
m17934 VDDREF 2325 2281 VDDREF pch l=0.04u w=0.8u
m17935 VDDREF 2347 2282 VDDREF pch l=0.04u w=0.8u
m17936 1931 2440 VDDREF VDDREF pch l=0.04u w=0.8u
m17937 VDDREF 2348 2283 VDDREF pch l=0.04u w=0.8u
m17938 VDDREF FBDIV[7] 2284 VDDREF pch l=0.04u w=0.8u
m17939 VDDREF 1876 2286 VDDREF pch l=0.04u w=0.8u
m17940 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m17941 2291 2192 2268 VDDREF pch l=0.04u w=0.8u
m17942 2292 2193 2269 VDDREF pch l=0.04u w=0.8u
m17943 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m17944 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m17945 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m17946 2293 292 VDDREF VDDREF pch l=0.04u w=0.8u
m17947 VDDREF 2326 1919 VDDREF pch l=0.04u w=0.8u
m17948 2294 1027 VDDREF VDDREF pch l=0.04u w=0.8u
m17949 VDDREF 2328 1921 VDDREF pch l=0.04u w=0.8u
m17950 VDDREF 2330 1923 VDDREF pch l=0.04u w=0.8u
m17951 VDDREF 2335 1927 VDDREF pch l=0.04u w=0.8u
m17952 VDDREF 2339 1931 VDDREF pch l=0.04u w=0.8u
m17953 2295 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17954 VDDREF 3736 2290 VDDREF pch l=0.04u w=0.8u
m17955 VDDREF 2400 VDDREF VDDREF pch l=0.26u w=1u
m17956 VDDREF 2401 VDDREF VDDREF pch l=0.26u w=1u
m17957 30174 4328 2291 VDDREF pch l=0.04u w=0.12u
m17958 30175 4328 2292 VDDREF pch l=0.04u w=0.12u
m17959 2296 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17960 2297 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17961 2298 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17962 2299 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m17963 2300 2270 VDDREF VDDREF pch l=0.04u w=0.8u
m17964 2301 2271 VDDREF VDDREF pch l=0.04u w=0.8u
m17965 2086 2486 VDDREF VDDREF pch l=0.04u w=0.8u
m17966 2289 2369 VDDREF VDDREF pch l=0.04u w=0.8u
m17967 2308 2342 VDDREF VDDREF pch l=0.04u w=0.8u
m17968 2309 2343 VDDREF VDDREF pch l=0.04u w=0.8u
m17969 2310 2274 VDDREF VDDREF pch l=0.04u w=0.8u
m17970 2311 2275 VDDREF VDDREF pch l=0.04u w=0.8u
m17971 2312 2276 VDDREF VDDREF pch l=0.04u w=0.8u
m17972 2313 2344 VDDREF VDDREF pch l=0.04u w=0.8u
m17973 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m17974 2314 131 VDDREF VDDREF pch l=0.04u w=0.8u
m17975 2315 2345 VDDREF VDDREF pch l=0.04u w=0.8u
m17976 2316 2346 VDDREF VDDREF pch l=0.04u w=0.8u
m17977 2317 2325 VDDREF VDDREF pch l=0.04u w=0.8u
m17978 2318 2347 VDDREF VDDREF pch l=0.04u w=0.8u
m17979 2319 2348 VDDREF VDDREF pch l=0.04u w=0.8u
m17980 2320 FBDIV[7] VDDREF VDDREF pch l=0.04u w=0.8u
m17981 VDDREF 2349 30174 VDDREF pch l=0.04u w=0.12u
m17982 VDDREF 2350 30175 VDDREF pch l=0.04u w=0.12u
m17983 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m17984 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m17985 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m17986 VDDREF 2304 2305 VDDREF pch l=0.04u w=1u
m17987 VDDREF 2307 2306 VDDREF pch l=0.04u w=1u
m17988 VDDREF 2648 2289 VDDREF pch l=0.04u w=0.8u
m17989 2302 110 292 VDDREF pch l=0.04u w=0.8u
m17990 2326 2198 VDDREF VDDREF pch l=0.04u w=0.8u
m17991 2303 2290 1027 VDDREF pch l=0.04u w=0.8u
m17992 2328 2200 VDDREF VDDREF pch l=0.04u w=0.8u
m17993 2330 2202 VDDREF VDDREF pch l=0.04u w=0.8u
m17994 2335 2206 VDDREF VDDREF pch l=0.04u w=0.8u
m17995 2339 2210 VDDREF VDDREF pch l=0.04u w=0.8u
m17996 2332 4328 2321 VDDREF pch l=0.04u w=0.8u
m17997 VDDREF 2400 VDDREF VDDREF pch l=0.26u w=1u
m17998 VDDREF 2401 VDDREF VDDREF pch l=0.26u w=1u
m17999 2349 2291 VDDREF VDDREF pch l=0.04u w=0.8u
m18000 2350 2292 VDDREF VDDREF pch l=0.04u w=0.8u
m18001 2351 4328 2322 VDDREF pch l=0.04u w=0.8u
m18002 2352 4328 2323 VDDREF pch l=0.04u w=0.8u
m18003 2353 4328 2324 VDDREF pch l=0.04u w=0.8u
m18004 2354 4328 2325 VDDREF pch l=0.04u w=0.8u
m18005 2355 2556 VDDREF VDDREF pch l=0.04u w=0.8u
m18006 2356 2557 VDDREF VDDREF pch l=0.04u w=0.8u
m18007 2357 2222 VDDREF VDDREF pch l=0.04u w=0.8u
m18008 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m18009 30197 2289 VDDREF VDDREF pch l=0.04u w=0.12u
m18010 110 292 2302 VDDREF pch l=0.04u w=0.8u
m18011 VDDREF 2239 2326 VDDREF pch l=0.04u w=0.8u
m18012 2290 1027 2303 VDDREF pch l=0.04u w=0.8u
m18013 VDDREF 2240 2328 VDDREF pch l=0.04u w=0.8u
m18014 VDDREF 2241 2330 VDDREF pch l=0.04u w=0.8u
m18015 VDDREF 2242 2335 VDDREF pch l=0.04u w=0.8u
m18016 VDDREF 2243 2339 VDDREF pch l=0.04u w=0.8u
m18017 2361 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18018 2362 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18019 2363 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18020 2327 2344 2342 VDDREF pch l=0.04u w=0.8u
m18021 2329 2357 2343 VDDREF pch l=0.04u w=0.8u
m18022 2364 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18023 2365 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18024 2366 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18025 2331 FRAC[7] 2344 VDDREF pch l=0.04u w=0.8u
m18026 30198 2295 2332 VDDREF pch l=0.04u w=0.12u
m18027 2333 2345 131 VDDREF pch l=0.04u w=0.8u
m18028 2334 2359 2345 VDDREF pch l=0.04u w=0.8u
m18029 2336 2324 2346 VDDREF pch l=0.04u w=0.8u
m18030 2337 2267 2325 VDDREF pch l=0.04u w=0.8u
m18031 2338 2360 2347 VDDREF pch l=0.04u w=0.8u
m18032 2340 FRAC[7] 2348 VDDREF pch l=0.04u w=0.8u
m18033 2341 2267 FBDIV[7] VDDREF pch l=0.04u w=0.8u
m18034 30201 2296 2351 VDDREF pch l=0.04u w=0.12u
m18035 30202 2297 2352 VDDREF pch l=0.04u w=0.12u
m18036 30203 2298 2353 VDDREF pch l=0.04u w=0.12u
m18037 30204 2299 2354 VDDREF pch l=0.04u w=0.12u
m18038 VDDREF 3012 2355 VDDREF pch l=0.04u w=0.8u
m18039 VDDREF 303 2356 VDDREF pch l=0.04u w=0.8u
m18040 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m18041 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m18042 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m18043 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18044 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18045 2369 2403 30197 VDDREF pch l=0.04u w=0.12u
m18046 VDDREF 2400 VDDREF VDDREF pch l=0.26u w=1u
m18047 VDDREF 2401 VDDREF VDDREF pch l=0.26u w=1u
m18048 2344 2342 2327 VDDREF pch l=0.04u w=0.8u
m18049 2357 2343 2329 VDDREF pch l=0.04u w=0.8u
m18050 FRAC[7] 2344 2331 VDDREF pch l=0.04u w=0.8u
m18051 VDDREF 2381 30198 VDDREF pch l=0.04u w=0.12u
m18052 2345 131 2333 VDDREF pch l=0.04u w=0.8u
m18053 2359 2345 2334 VDDREF pch l=0.04u w=0.8u
m18054 2324 2346 2336 VDDREF pch l=0.04u w=0.8u
m18055 2267 2325 2337 VDDREF pch l=0.04u w=0.8u
m18056 2360 2347 2338 VDDREF pch l=0.04u w=0.8u
m18057 FRAC[7] 2348 2340 VDDREF pch l=0.04u w=0.8u
m18058 2267 FBDIV[7] 2341 VDDREF pch l=0.04u w=0.8u
m18059 VDDREF 2349 2367 VDDREF pch l=0.04u w=0.8u
m18060 VDDREF 2350 2368 VDDREF pch l=0.04u w=0.8u
m18061 VDDREF 2392 30201 VDDREF pch l=0.04u w=0.12u
m18062 VDDREF 2393 30202 VDDREF pch l=0.04u w=0.12u
m18063 VDDREF 2394 30203 VDDREF pch l=0.04u w=0.12u
m18064 VDDREF 2395 30204 VDDREF pch l=0.04u w=0.12u
m18065 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m18066 2188 2454 2369 VDDREF pch l=0.04u w=0.8u
m18067 2370 2302 VDDREF VDDREF pch l=0.04u w=0.8u
m18068 2239 395 2222 VDDREF pch l=0.04u w=0.8u
m18069 2371 2303 VDDREF VDDREF pch l=0.04u w=0.8u
m18070 2240 2225 139 VDDREF pch l=0.04u w=0.8u
m18071 2241 2222 FRAC[17] VDDREF pch l=0.04u w=0.8u
m18072 2381 2332 VDDREF VDDREF pch l=0.04u w=0.8u
m18073 2242 1941 1815 VDDREF pch l=0.04u w=0.8u
m18074 2243 1942 FRAC[17] VDDREF pch l=0.04u w=0.8u
m18075 2375 4328 2373 VDDREF pch l=0.04u w=0.8u
m18076 2376 4328 2374 VDDREF pch l=0.04u w=0.8u
m18077 2377 4328 296 VDDREF pch l=0.04u w=0.8u
m18078 2378 4328 2310 VDDREF pch l=0.04u w=0.8u
m18079 2379 4328 2311 VDDREF pch l=0.04u w=0.8u
m18080 2380 4328 2312 VDDREF pch l=0.04u w=0.8u
m18081 710 2367 VDDREF VDDREF pch l=0.04u w=0.8u
m18082 1086 2368 VDDREF VDDREF pch l=0.04u w=0.8u
m18083 2392 2351 VDDREF VDDREF pch l=0.04u w=0.8u
m18084 2393 2352 VDDREF VDDREF pch l=0.04u w=0.8u
m18085 2394 2353 VDDREF VDDREF pch l=0.04u w=0.8u
m18086 2395 2354 VDDREF VDDREF pch l=0.04u w=0.8u
m18087 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m18088 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m18089 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m18090 2396 2300 VDDREF VDDREF pch l=0.04u w=0.8u
m18091 2397 2301 VDDREF VDDREF pch l=0.04u w=0.8u
m18092 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18093 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18094 VDDREF 2400 VDDREF VDDREF pch l=0.26u w=1u
m18095 VDDREF 2401 VDDREF VDDREF pch l=0.26u w=1u
m18096 VDDREF 2143 2370 VDDREF pch l=0.04u w=0.8u
m18097 395 2222 2239 VDDREF pch l=0.04u w=0.8u
m18098 VDDREF 2147 2371 VDDREF pch l=0.04u w=0.8u
m18099 2225 139 2240 VDDREF pch l=0.04u w=0.8u
m18100 2222 FRAC[17] 2241 VDDREF pch l=0.04u w=0.8u
m18101 1941 1815 2242 VDDREF pch l=0.04u w=0.8u
m18102 1942 FRAC[17] 2243 VDDREF pch l=0.04u w=0.8u
m18103 30221 2361 2375 VDDREF pch l=0.04u w=0.12u
m18104 30222 2362 2376 VDDREF pch l=0.04u w=0.12u
m18105 30223 2363 2377 VDDREF pch l=0.04u w=0.12u
m18106 2382 2327 VDDREF VDDREF pch l=0.04u w=0.8u
m18107 2383 2329 VDDREF VDDREF pch l=0.04u w=0.8u
m18108 30224 2364 2378 VDDREF pch l=0.04u w=0.12u
m18109 30225 2365 2379 VDDREF pch l=0.04u w=0.12u
m18110 30226 2366 2380 VDDREF pch l=0.04u w=0.12u
m18111 2384 2331 VDDREF VDDREF pch l=0.04u w=0.8u
m18112 2385 2333 VDDREF VDDREF pch l=0.04u w=0.8u
m18113 2386 2334 VDDREF VDDREF pch l=0.04u w=0.8u
m18114 2387 2336 VDDREF VDDREF pch l=0.04u w=0.8u
m18115 2388 2337 VDDREF VDDREF pch l=0.04u w=0.8u
m18116 2389 2338 VDDREF VDDREF pch l=0.04u w=0.8u
m18117 2390 2340 VDDREF VDDREF pch l=0.04u w=0.8u
m18118 2391 2341 VDDREF VDDREF pch l=0.04u w=0.8u
m18119 2398 155 VDDREF VDDREF pch l=0.04u w=0.8u
m18120 VDDREF 2300 2396 VDDREF pch l=0.04u w=0.8u
m18121 VDDREF 2301 2397 VDDREF pch l=0.04u w=0.8u
m18122 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m18123 2399 2399 VDDREF VDDREF pch l=0.04u w=1u
m18124 2402 2402 VDDREF VDDREF pch l=0.04u w=1u
m18125 2403 2454 VDDREF VDDREF pch l=0.04u w=0.8u
m18126 VDDREF 2418 30221 VDDREF pch l=0.04u w=0.12u
m18127 VDDREF 2419 30222 VDDREF pch l=0.04u w=0.12u
m18128 VDDREF 2420 30223 VDDREF pch l=0.04u w=0.12u
m18129 VDDREF 2159 2382 VDDREF pch l=0.04u w=0.8u
m18130 VDDREF 2161 2383 VDDREF pch l=0.04u w=0.8u
m18131 VDDREF 2422 30224 VDDREF pch l=0.04u w=0.12u
m18132 VDDREF 2423 30225 VDDREF pch l=0.04u w=0.12u
m18133 VDDREF 2424 30226 VDDREF pch l=0.04u w=0.12u
m18134 VDDREF 2163 2384 VDDREF pch l=0.04u w=0.8u
m18135 2404 2295 2381 VDDREF pch l=0.04u w=0.8u
m18136 VDDREF 2164 2385 VDDREF pch l=0.04u w=0.8u
m18137 VDDREF 2165 2386 VDDREF pch l=0.04u w=0.8u
m18138 VDDREF 2167 2387 VDDREF pch l=0.04u w=0.8u
m18139 VDDREF 2168 2388 VDDREF pch l=0.04u w=0.8u
m18140 VDDREF 2169 2389 VDDREF pch l=0.04u w=0.8u
m18141 VDDREF 2171 2390 VDDREF pch l=0.04u w=0.8u
m18142 VDDREF 2172 2391 VDDREF pch l=0.04u w=0.8u
m18143 2410 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18144 2411 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18145 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m18146 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m18147 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m18148 2412 2296 2392 VDDREF pch l=0.04u w=0.8u
m18149 2413 2297 2393 VDDREF pch l=0.04u w=0.8u
m18150 2414 2298 2394 VDDREF pch l=0.04u w=0.8u
m18151 2415 2299 2395 VDDREF pch l=0.04u w=0.8u
m18152 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18153 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18154 2417 2370 VDDREF VDDREF pch l=0.04u w=0.8u
m18155 2418 2375 VDDREF VDDREF pch l=0.04u w=0.8u
m18156 2419 2376 VDDREF VDDREF pch l=0.04u w=0.8u
m18157 2420 2377 VDDREF VDDREF pch l=0.04u w=0.8u
m18158 VDDREF 395 2405 VDDREF pch l=0.04u w=0.8u
m18159 2421 2371 VDDREF VDDREF pch l=0.04u w=0.8u
m18160 VDDREF 2225 2406 VDDREF pch l=0.04u w=0.8u
m18161 2422 2378 VDDREF VDDREF pch l=0.04u w=0.8u
m18162 2423 2379 VDDREF VDDREF pch l=0.04u w=0.8u
m18163 2424 2380 VDDREF VDDREF pch l=0.04u w=0.8u
m18164 VDDREF 2222 2407 VDDREF pch l=0.04u w=0.8u
m18165 30243 4328 2404 VDDREF pch l=0.04u w=0.12u
m18166 VDDREF 1941 2408 VDDREF pch l=0.04u w=0.8u
m18167 VDDREF 1942 2409 VDDREF pch l=0.04u w=0.8u
m18168 2425 155 VDDREF VDDREF pch l=0.04u w=0.8u
m18169 30250 4328 2412 VDDREF pch l=0.04u w=0.12u
m18170 30251 4328 2413 VDDREF pch l=0.04u w=0.12u
m18171 30252 4328 2414 VDDREF pch l=0.04u w=0.12u
m18172 30253 4328 2415 VDDREF pch l=0.04u w=0.12u
m18173 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m18174 2426 2396 VDDREF VDDREF pch l=0.04u w=0.8u
m18175 2427 2397 VDDREF VDDREF pch l=0.04u w=0.8u
m18176 VDDREF 2454 2416 VDDREF pch l=0.04u w=0.8u
m18177 VDDREF 2261 2417 VDDREF pch l=0.04u w=0.8u
m18178 VDDREF 2262 2421 VDDREF pch l=0.04u w=0.8u
m18179 VDDREF 2453 30243 VDDREF pch l=0.04u w=0.12u
m18180 2429 2382 VDDREF VDDREF pch l=0.04u w=0.8u
m18181 2431 2383 VDDREF VDDREF pch l=0.04u w=0.8u
m18182 2433 2384 VDDREF VDDREF pch l=0.04u w=0.8u
m18183 2434 2385 VDDREF VDDREF pch l=0.04u w=0.8u
m18184 2435 2386 VDDREF VDDREF pch l=0.04u w=0.8u
m18185 2437 2387 VDDREF VDDREF pch l=0.04u w=0.8u
m18186 2438 2388 VDDREF VDDREF pch l=0.04u w=0.8u
m18187 2439 2389 VDDREF VDDREF pch l=0.04u w=0.8u
m18188 2441 2390 VDDREF VDDREF pch l=0.04u w=0.8u
m18189 2442 2391 VDDREF VDDREF pch l=0.04u w=0.8u
m18190 VDDREF FBDIV[7] 2425 VDDREF pch l=0.04u w=0.8u
m18191 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m18192 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m18193 VDDREF 2455 VDDREF VDDREF pch l=0.26u w=1u
m18194 2443 4328 2349 VDDREF pch l=0.04u w=0.8u
m18195 2444 4328 2350 VDDREF pch l=0.04u w=0.8u
m18196 VDDREF 2346 30250 VDDREF pch l=0.04u w=0.12u
m18197 VDDREF 2345 30251 VDDREF pch l=0.04u w=0.12u
m18198 VDDREF 2348 30252 VDDREF pch l=0.04u w=0.12u
m18199 VDDREF 2347 30253 VDDREF pch l=0.04u w=0.12u
m18200 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18201 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18202 VDDREF 2396 2426 VDDREF pch l=0.04u w=0.8u
m18203 VDDREF 2397 2427 VDDREF pch l=0.04u w=0.8u
m18204 2445 3454 VDDREF VDDREF pch l=0.04u w=0.8u
m18205 2446 2508 VDDREF VDDREF pch l=0.04u w=0.8u
m18206 2453 2404 VDDREF VDDREF pch l=0.04u w=0.8u
m18207 2447 2361 2418 VDDREF pch l=0.04u w=0.8u
m18208 2448 2362 2419 VDDREF pch l=0.04u w=0.8u
m18209 2449 2363 2420 VDDREF pch l=0.04u w=0.8u
m18210 2428 395 VDDREF VDDREF pch l=0.04u w=0.8u
m18211 VDDREF 2272 2429 VDDREF pch l=0.04u w=0.8u
m18212 2430 2225 VDDREF VDDREF pch l=0.04u w=0.8u
m18213 VDDREF 2273 2431 VDDREF pch l=0.04u w=0.8u
m18214 2450 2364 2422 VDDREF pch l=0.04u w=0.8u
m18215 2451 2365 2423 VDDREF pch l=0.04u w=0.8u
m18216 2452 2366 2424 VDDREF pch l=0.04u w=0.8u
m18217 2432 2222 VDDREF VDDREF pch l=0.04u w=0.8u
m18218 VDDREF 2277 2433 VDDREF pch l=0.04u w=0.8u
m18219 VDDREF 2278 2434 VDDREF pch l=0.04u w=0.8u
m18220 VDDREF 2279 2435 VDDREF pch l=0.04u w=0.8u
m18221 2436 1941 VDDREF VDDREF pch l=0.04u w=0.8u
m18222 VDDREF 2280 2437 VDDREF pch l=0.04u w=0.8u
m18223 VDDREF 2281 2438 VDDREF pch l=0.04u w=0.8u
m18224 VDDREF 2282 2439 VDDREF pch l=0.04u w=0.8u
m18225 2440 1942 VDDREF VDDREF pch l=0.04u w=0.8u
m18226 VDDREF 2283 2441 VDDREF pch l=0.04u w=0.8u
m18227 VDDREF 2284 2442 VDDREF pch l=0.04u w=0.8u
m18228 2456 2456 VDDREF VDDREF pch l=0.04u w=1u
m18229 30261 2410 2443 VDDREF pch l=0.04u w=0.12u
m18230 30262 2411 2444 VDDREF pch l=0.04u w=0.12u
m18231 VDDREF 2463 VDDREF VDDREF pch l=0.26u w=1u
m18232 2346 2412 VDDREF VDDREF pch l=0.04u w=0.8u
m18233 2345 2413 VDDREF VDDREF pch l=0.04u w=0.8u
m18234 2348 2414 VDDREF VDDREF pch l=0.04u w=0.8u
m18235 2347 2415 VDDREF VDDREF pch l=0.04u w=0.8u
m18236 2426 2396 VDDREF VDDREF pch l=0.04u w=0.8u
m18237 2427 2397 VDDREF VDDREF pch l=0.04u w=0.8u
m18238 VDDREF 1918 2446 VDDREF pch l=0.04u w=0.8u
m18239 2454 2487 VDDREF VDDREF pch l=0.04u w=0.8u
m18240 2457 2302 VDDREF VDDREF pch l=0.04u w=0.8u
m18241 30270 4328 2447 VDDREF pch l=0.04u w=0.12u
m18242 30271 4328 2448 VDDREF pch l=0.04u w=0.12u
m18243 30272 4328 2449 VDDREF pch l=0.04u w=0.12u
m18244 VDDREF 2222 2428 VDDREF pch l=0.04u w=0.8u
m18245 2458 2303 VDDREF VDDREF pch l=0.04u w=0.8u
m18246 VDDREF 139 2430 VDDREF pch l=0.04u w=0.8u
m18247 30273 4328 2450 VDDREF pch l=0.04u w=0.12u
m18248 30274 4328 2451 VDDREF pch l=0.04u w=0.12u
m18249 30275 4328 2452 VDDREF pch l=0.04u w=0.12u
m18250 VDDREF FRAC[17] 2432 VDDREF pch l=0.04u w=0.8u
m18251 VDDREF 1815 2436 VDDREF pch l=0.04u w=0.8u
m18252 VDDREF FRAC[17] 2440 VDDREF pch l=0.04u w=0.8u
m18253 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m18254 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m18255 2459 2398 VDDREF VDDREF pch l=0.04u w=0.8u
m18256 VDDREF 2481 30261 VDDREF pch l=0.04u w=0.12u
m18257 VDDREF 2482 30262 VDDREF pch l=0.04u w=0.12u
m18258 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18259 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18260 2462 2462 VDDREF VDDREF pch l=0.04u w=1u
m18261 VDDREF 2396 2426 VDDREF pch l=0.04u w=0.8u
m18262 VDDREF 2397 2427 VDDREF pch l=0.04u w=0.8u
m18263 VDDREF 2648 2454 VDDREF pch l=0.04u w=0.8u
m18264 2464 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m18265 VDDREF 91 30270 VDDREF pch l=0.04u w=0.12u
m18266 VDDREF 2342 30271 VDDREF pch l=0.04u w=0.12u
m18267 VDDREF 125 30272 VDDREF pch l=0.04u w=0.12u
m18268 VDDREF 2486 30273 VDDREF pch l=0.04u w=0.12u
m18269 VDDREF 2344 30274 VDDREF pch l=0.04u w=0.12u
m18270 VDDREF 129 30275 VDDREF pch l=0.04u w=0.12u
m18271 2467 2327 VDDREF VDDREF pch l=0.04u w=0.8u
m18272 2469 2329 VDDREF VDDREF pch l=0.04u w=0.8u
m18273 2471 2331 VDDREF VDDREF pch l=0.04u w=0.8u
m18274 2472 2333 VDDREF VDDREF pch l=0.04u w=0.8u
m18275 2473 2334 VDDREF VDDREF pch l=0.04u w=0.8u
m18276 2475 2336 VDDREF VDDREF pch l=0.04u w=0.8u
m18277 2476 2337 VDDREF VDDREF pch l=0.04u w=0.8u
m18278 2477 2338 VDDREF VDDREF pch l=0.04u w=0.8u
m18279 2479 2340 VDDREF VDDREF pch l=0.04u w=0.8u
m18280 2480 2341 VDDREF VDDREF pch l=0.04u w=0.8u
m18281 VDDREF 2453 2459 VDDREF pch l=0.04u w=0.8u
m18282 2481 2443 VDDREF VDDREF pch l=0.04u w=0.8u
m18283 2482 2444 VDDREF VDDREF pch l=0.04u w=0.8u
m18284 VDDREF 2460 2461 VDDREF pch l=0.04u w=1u
m18285 2426 2396 VDDREF VDDREF pch l=0.04u w=0.8u
m18286 2427 2397 VDDREF VDDREF pch l=0.04u w=0.8u
m18287 VDDREF 1918 2464 VDDREF pch l=0.04u w=0.8u
m18288 2485 1918 VDDREF VDDREF pch l=0.04u w=0.8u
m18289 91 2447 VDDREF VDDREF pch l=0.04u w=0.8u
m18290 2342 2448 VDDREF VDDREF pch l=0.04u w=0.8u
m18291 VDDREF 2492 VDDREF VDDREF pch l=0.26u w=1u
m18292 125 2449 VDDREF VDDREF pch l=0.04u w=0.8u
m18293 2486 2450 VDDREF VDDREF pch l=0.04u w=0.8u
m18294 2344 2451 VDDREF VDDREF pch l=0.04u w=0.8u
m18295 VDDREF 2494 VDDREF VDDREF pch l=0.26u w=1u
m18296 129 2452 VDDREF VDDREF pch l=0.04u w=0.8u
m18297 2465 2143 2302 VDDREF pch l=0.04u w=0.8u
m18298 2373 2496 2466 VDDREF pch l=0.04u w=0.8u
m18299 1041 2147 2303 VDDREF pch l=0.04u w=0.8u
m18300 2488 2497 2468 VDDREF pch l=0.04u w=0.8u
m18301 2490 2498 2470 VDDREF pch l=0.04u w=0.8u
m18302 2153 2499 2474 VDDREF pch l=0.04u w=0.8u
m18303 2155 2500 2478 VDDREF pch l=0.04u w=0.8u
m18304 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18305 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18306 VDDREF 2484 2483 VDDREF pch l=0.04u w=1u
m18307 VDDREF 2396 2426 VDDREF pch l=0.04u w=0.8u
m18308 VDDREF 2397 2427 VDDREF pch l=0.04u w=0.8u
m18309 2493 2493 VDDREF VDDREF pch l=0.04u w=1u
m18310 2495 2495 VDDREF VDDREF pch l=0.04u w=1u
m18311 VDDREF 2524 2487 VDDREF pch l=0.04u w=0.8u
m18312 2143 2302 2465 VDDREF pch l=0.04u w=0.8u
m18313 2496 2466 2373 VDDREF pch l=0.04u w=0.8u
m18314 2147 2303 1041 VDDREF pch l=0.04u w=0.8u
m18315 2497 2468 2488 VDDREF pch l=0.04u w=0.8u
m18316 2498 2470 2490 VDDREF pch l=0.04u w=0.8u
m18317 2499 2474 2153 VDDREF pch l=0.04u w=0.8u
m18318 2500 2478 2155 VDDREF pch l=0.04u w=0.8u
m18319 2374 2159 2327 VDDREF pch l=0.04u w=0.8u
m18320 2489 2161 2329 VDDREF pch l=0.04u w=0.8u
m18321 2343 2163 2331 VDDREF pch l=0.04u w=0.8u
m18322 2321 2164 2333 VDDREF pch l=0.04u w=0.8u
m18323 2323 2165 2334 VDDREF pch l=0.04u w=0.8u
m18324 2322 2167 2336 VDDREF pch l=0.04u w=0.8u
m18325 2359 2168 2337 VDDREF pch l=0.04u w=0.8u
m18326 2325 2169 2338 VDDREF pch l=0.04u w=0.8u
m18327 2324 2171 2340 VDDREF pch l=0.04u w=0.8u
m18328 2360 2172 2341 VDDREF pch l=0.04u w=0.8u
m18329 2501 2459 VDDREF VDDREF pch l=0.04u w=0.8u
m18330 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18331 2504 2410 2481 VDDREF pch l=0.04u w=0.8u
m18332 2505 2411 2482 VDDREF pch l=0.04u w=0.8u
m18333 2426 2396 VDDREF VDDREF pch l=0.04u w=0.8u
m18334 2427 2397 VDDREF VDDREF pch l=0.04u w=0.8u
m18335 30313 2416 VDDREF VDDREF pch l=0.04u w=0.24u
m18336 2509 2464 VDDREF VDDREF pch l=0.04u w=0.8u
m18337 2491 2508 1918 VDDREF pch l=0.04u w=0.8u
m18338 2510 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18339 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18340 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18341 2159 2327 2374 VDDREF pch l=0.04u w=0.8u
m18342 2161 2329 2489 VDDREF pch l=0.04u w=0.8u
m18343 2163 2331 2343 VDDREF pch l=0.04u w=0.8u
m18344 2164 2333 2321 VDDREF pch l=0.04u w=0.8u
m18345 2165 2334 2323 VDDREF pch l=0.04u w=0.8u
m18346 2167 2336 2322 VDDREF pch l=0.04u w=0.8u
m18347 2168 2337 2359 VDDREF pch l=0.04u w=0.8u
m18348 2169 2338 2325 VDDREF pch l=0.04u w=0.8u
m18349 2171 2340 2324 VDDREF pch l=0.04u w=0.8u
m18350 2172 2341 2360 VDDREF pch l=0.04u w=0.8u
m18351 VDDREF 2425 2501 VDDREF pch l=0.04u w=0.8u
m18352 VDDREF 2503 2502 VDDREF pch l=0.04u w=1u
m18353 30318 4328 2504 VDDREF pch l=0.04u w=0.12u
m18354 30319 4328 2505 VDDREF pch l=0.04u w=0.12u
m18355 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18356 VDDREF 2396 2426 VDDREF pch l=0.04u w=0.8u
m18357 VDDREF 2397 2427 VDDREF pch l=0.04u w=0.8u
m18358 VDDREF 2506 2507 VDDREF pch l=0.04u w=1u
m18359 2524 5232 30313 VDDREF pch l=0.04u w=0.24u
m18360 2508 1918 2491 VDDREF pch l=0.04u w=0.8u
m18361 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18362 2525 2417 VDDREF VDDREF pch l=0.04u w=0.8u
m18363 VDDREF 2496 2511 VDDREF pch l=0.04u w=0.8u
m18364 2526 2421 VDDREF VDDREF pch l=0.04u w=0.8u
m18365 VDDREF 2497 2512 VDDREF pch l=0.04u w=0.8u
m18366 VDDREF 2498 2513 VDDREF pch l=0.04u w=0.8u
m18367 VDDREF 2515 2514 VDDREF pch l=0.04u w=1u
m18368 VDDREF 2516 2517 VDDREF pch l=0.04u w=1u
m18369 VDDREF 2499 2518 VDDREF pch l=0.04u w=0.8u
m18370 VDDREF 2520 2519 VDDREF pch l=0.04u w=1u
m18371 VDDREF 2521 2522 VDDREF pch l=0.04u w=1u
m18372 VDDREF 2500 2523 VDDREF pch l=0.04u w=0.8u
m18373 VDDREF 2554 30318 VDDREF pch l=0.04u w=0.12u
m18374 VDDREF 2555 30319 VDDREF pch l=0.04u w=0.12u
m18375 VDDREF 2558 VDDREF VDDREF pch l=0.26u w=1u
m18376 VDDREF 2561 VDDREF VDDREF pch l=0.26u w=1u
m18377 2541 2615 2524 VDDREF pch l=0.04u w=0.8u
m18378 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18379 2542 4328 LOCK VDDREF pch l=0.04u w=0.8u
m18380 2544 2429 VDDREF VDDREF pch l=0.04u w=0.8u
m18381 2545 2431 VDDREF VDDREF pch l=0.04u w=0.8u
m18382 2546 2433 VDDREF VDDREF pch l=0.04u w=0.8u
m18383 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18384 2547 2434 VDDREF VDDREF pch l=0.04u w=0.8u
m18385 2548 2435 VDDREF VDDREF pch l=0.04u w=0.8u
m18386 2549 2437 VDDREF VDDREF pch l=0.04u w=0.8u
m18387 2550 2438 VDDREF VDDREF pch l=0.04u w=0.8u
m18388 2551 2439 VDDREF VDDREF pch l=0.04u w=0.8u
m18389 2552 2441 VDDREF VDDREF pch l=0.04u w=0.8u
m18390 2553 2442 VDDREF VDDREF pch l=0.04u w=0.8u
m18391 2554 2504 VDDREF VDDREF pch l=0.04u w=0.8u
m18392 2555 2505 VDDREF VDDREF pch l=0.04u w=0.8u
m18393 VDDREF 2527 2528 VDDREF pch l=0.04u w=1u
m18394 VDDREF 2530 2529 VDDREF pch l=0.04u w=1u
m18395 VDDREF 2531 2532 VDDREF pch l=0.04u w=1u
m18396 VDDREF 2534 2533 VDDREF pch l=0.04u w=1u
m18397 VDDREF 2535 2536 VDDREF pch l=0.04u w=1u
m18398 VDDREF 2538 2537 VDDREF pch l=0.04u w=1u
m18399 VDDREF 2539 2540 VDDREF pch l=0.04u w=1u
m18400 2556 2716 VDDREF VDDREF pch l=0.04u w=0.8u
m18401 2557 2716 VDDREF VDDREF pch l=0.04u w=0.8u
m18402 VDDREF 2631 VDDREF VDDREF pch l=0.26u w=1u
m18403 2559 2559 VDDREF VDDREF pch l=0.04u w=1u
m18404 2560 2560 VDDREF VDDREF pch l=0.04u w=1u
m18405 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18406 VDDREF 2641 VDDREF VDDREF pch l=0.26u w=1u
m18407 VDDREF 2642 VDDREF VDDREF pch l=0.26u w=1u
m18408 VDDREF 2645 VDDREF VDDREF pch l=0.26u w=1u
m18409 VDDREF 2646 VDDREF VDDREF pch l=0.26u w=1u
m18410 2543 2491 VDDREF VDDREF pch l=0.04u w=0.8u
m18411 30336 2510 2542 VDDREF pch l=0.04u w=0.12u
m18412 2562 1464 VDDREF VDDREF pch l=0.04u w=0.8u
m18413 2198 2669 VDDREF VDDREF pch l=0.04u w=0.8u
m18414 2563 1465 VDDREF VDDREF pch l=0.04u w=0.8u
m18415 2200 2670 VDDREF VDDREF pch l=0.04u w=0.8u
m18416 2202 2671 VDDREF VDDREF pch l=0.04u w=0.8u
m18417 2206 2672 VDDREF VDDREF pch l=0.04u w=0.8u
m18418 2210 2673 VDDREF VDDREF pch l=0.04u w=0.8u
m18419 VDDREF 2270 2556 VDDREF pch l=0.04u w=0.8u
m18420 VDDREF 2271 2557 VDDREF pch l=0.04u w=0.8u
m18421 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18422 2541 2594 VDDREF VDDREF pch l=0.04u w=0.8u
m18423 VDDREF 2630 2543 VDDREF pch l=0.04u w=0.8u
m18424 VDDREF 2580 30336 VDDREF pch l=0.04u w=0.12u
m18425 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18426 VDDREF 1755 2562 VDDREF pch l=0.04u w=0.8u
m18427 VDDREF 2584 2198 VDDREF pch l=0.04u w=0.8u
m18428 VDDREF 1756 2563 VDDREF pch l=0.04u w=0.8u
m18429 VDDREF 2585 2200 VDDREF pch l=0.04u w=0.8u
m18430 VDDREF 2586 2202 VDDREF pch l=0.04u w=0.8u
m18431 VDDREF 2587 2206 VDDREF pch l=0.04u w=0.8u
m18432 VDDREF 2588 2210 VDDREF pch l=0.04u w=0.8u
m18433 2568 1488 VDDREF VDDREF pch l=0.04u w=0.8u
m18434 2569 1489 VDDREF VDDREF pch l=0.04u w=0.8u
m18435 2570 1490 VDDREF VDDREF pch l=0.04u w=0.8u
m18436 2571 1492 VDDREF VDDREF pch l=0.04u w=0.8u
m18437 2572 1493 VDDREF VDDREF pch l=0.04u w=0.8u
m18438 2573 1494 VDDREF VDDREF pch l=0.04u w=0.8u
m18439 2574 1495 VDDREF VDDREF pch l=0.04u w=0.8u
m18440 2575 1496 VDDREF VDDREF pch l=0.04u w=0.8u
m18441 2576 1497 VDDREF VDDREF pch l=0.04u w=0.8u
m18442 2577 1498 VDDREF VDDREF pch l=0.04u w=0.8u
m18443 2578 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18444 2579 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18445 VDDREF 2652 VDDREF VDDREF pch l=0.26u w=1u
m18446 VDDREF 2655 VDDREF VDDREF pch l=0.26u w=1u
m18447 VDDREF 2656 VDDREF VDDREF pch l=0.26u w=1u
m18448 VDDREF 2659 VDDREF VDDREF pch l=0.26u w=1u
m18449 VDDREF 2660 VDDREF VDDREF pch l=0.26u w=1u
m18450 VDDREF 2663 VDDREF VDDREF pch l=0.26u w=1u
m18451 VDDREF 2664 VDDREF VDDREF pch l=0.26u w=1u
m18452 VDDREF 2631 VDDREF VDDREF pch l=0.26u w=1u
m18453 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18454 VDDREF 2641 VDDREF VDDREF pch l=0.26u w=1u
m18455 VDDREF 2642 VDDREF VDDREF pch l=0.26u w=1u
m18456 VDDREF 2645 VDDREF VDDREF pch l=0.26u w=1u
m18457 VDDREF 2646 VDDREF VDDREF pch l=0.26u w=1u
m18458 VDDREF 2564 2565 VDDREF pch l=0.04u w=1u
m18459 VDDREF 2567 2566 VDDREF pch l=0.04u w=1u
m18460 VDDREF 2648 2541 VDDREF pch l=0.04u w=0.8u
m18461 2580 2542 VDDREF VDDREF pch l=0.04u w=0.8u
m18462 2562 2038 VDDREF VDDREF pch l=0.04u w=0.8u
m18463 2563 2039 VDDREF VDDREF pch l=0.04u w=0.8u
m18464 VDDREF 1774 2568 VDDREF pch l=0.04u w=0.8u
m18465 VDDREF 1776 2569 VDDREF pch l=0.04u w=0.8u
m18466 VDDREF 1778 2570 VDDREF pch l=0.04u w=0.8u
m18467 VDDREF 1780 2571 VDDREF pch l=0.04u w=0.8u
m18468 VDDREF 1781 2572 VDDREF pch l=0.04u w=0.8u
m18469 VDDREF 1783 2573 VDDREF pch l=0.04u w=0.8u
m18470 VDDREF 1784 2574 VDDREF pch l=0.04u w=0.8u
m18471 VDDREF 1785 2575 VDDREF pch l=0.04u w=0.8u
m18472 VDDREF 1787 2576 VDDREF pch l=0.04u w=0.8u
m18473 VDDREF 1788 2577 VDDREF pch l=0.04u w=0.8u
m18474 2581 4353 VDDREF VDDREF pch l=0.04u w=0.8u
m18475 2582 11 VDDREF VDDREF pch l=0.04u w=0.8u
m18476 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18477 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18478 30359 2541 VDDREF VDDREF pch l=0.04u w=0.12u
m18479 2583 2543 VDDREF VDDREF pch l=0.04u w=0.8u
m18480 2584 2466 VDDREF VDDREF pch l=0.04u w=0.8u
m18481 2568 2056 VDDREF VDDREF pch l=0.04u w=0.8u
m18482 2585 2468 VDDREF VDDREF pch l=0.04u w=0.8u
m18483 2569 2058 VDDREF VDDREF pch l=0.04u w=0.8u
m18484 2586 2470 VDDREF VDDREF pch l=0.04u w=0.8u
m18485 2570 2060 VDDREF VDDREF pch l=0.04u w=0.8u
m18486 2571 2062 VDDREF VDDREF pch l=0.04u w=0.8u
m18487 2572 2063 VDDREF VDDREF pch l=0.04u w=0.8u
m18488 2587 2474 VDDREF VDDREF pch l=0.04u w=0.8u
m18489 2573 2065 VDDREF VDDREF pch l=0.04u w=0.8u
m18490 2574 2066 VDDREF VDDREF pch l=0.04u w=0.8u
m18491 2575 2067 VDDREF VDDREF pch l=0.04u w=0.8u
m18492 2588 2478 VDDREF VDDREF pch l=0.04u w=0.8u
m18493 2576 2069 VDDREF VDDREF pch l=0.04u w=0.8u
m18494 2577 2070 VDDREF VDDREF pch l=0.04u w=0.8u
m18495 VDDREF 2652 VDDREF VDDREF pch l=0.26u w=1u
m18496 VDDREF 2655 VDDREF VDDREF pch l=0.26u w=1u
m18497 VDDREF 2656 VDDREF VDDREF pch l=0.26u w=1u
m18498 VDDREF 2659 VDDREF VDDREF pch l=0.26u w=1u
m18499 VDDREF 2660 VDDREF VDDREF pch l=0.26u w=1u
m18500 VDDREF 2663 VDDREF VDDREF pch l=0.26u w=1u
m18501 VDDREF 2664 VDDREF VDDREF pch l=0.26u w=1u
m18502 2589 4328 2554 VDDREF pch l=0.04u w=0.8u
m18503 2590 4328 2555 VDDREF pch l=0.04u w=0.8u
m18504 VDDREF 2631 VDDREF VDDREF pch l=0.26u w=1u
m18505 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18506 VDDREF 2641 VDDREF VDDREF pch l=0.26u w=1u
m18507 VDDREF 2642 VDDREF VDDREF pch l=0.26u w=1u
m18508 VDDREF 2645 VDDREF VDDREF pch l=0.26u w=1u
m18509 VDDREF 2646 VDDREF VDDREF pch l=0.26u w=1u
m18510 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18511 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18512 2594 2615 30359 VDDREF pch l=0.04u w=0.12u
m18513 VDDREF 2446 2583 VDDREF pch l=0.04u w=0.8u
m18514 2593 2510 2580 VDDREF pch l=0.04u w=0.8u
m18515 2595 2562 VDDREF VDDREF pch l=0.04u w=0.8u
m18516 VDDREF 2496 2584 VDDREF pch l=0.04u w=0.8u
m18517 2596 2563 VDDREF VDDREF pch l=0.04u w=0.8u
m18518 VDDREF 2497 2585 VDDREF pch l=0.04u w=0.8u
m18519 VDDREF 2498 2586 VDDREF pch l=0.04u w=0.8u
m18520 VDDREF 2499 2587 VDDREF pch l=0.04u w=0.8u
m18521 VDDREF 2500 2588 VDDREF pch l=0.04u w=0.8u
m18522 30371 2578 2589 VDDREF pch l=0.04u w=0.12u
m18523 30372 2579 2590 VDDREF pch l=0.04u w=0.12u
m18524 VDDREF 2592 2591 VDDREF pch l=0.04u w=1u
m18525 2597 4353 2355 VDDREF pch l=0.04u w=0.8u
m18526 2598 11 2356 VDDREF pch l=0.04u w=0.8u
m18527 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18528 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18529 2454 5232 2594 VDDREF pch l=0.04u w=0.8u
m18530 30375 4328 2593 VDDREF pch l=0.04u w=0.12u
m18531 VDDREF 2652 VDDREF VDDREF pch l=0.26u w=1u
m18532 VDDREF 2655 VDDREF VDDREF pch l=0.26u w=1u
m18533 VDDREF 2656 VDDREF VDDREF pch l=0.26u w=1u
m18534 VDDREF 2659 VDDREF VDDREF pch l=0.26u w=1u
m18535 VDDREF 2660 VDDREF VDDREF pch l=0.26u w=1u
m18536 VDDREF 2663 VDDREF VDDREF pch l=0.26u w=1u
m18537 VDDREF 2664 VDDREF VDDREF pch l=0.26u w=1u
m18538 2599 2568 VDDREF VDDREF pch l=0.04u w=0.8u
m18539 2600 2569 VDDREF VDDREF pch l=0.04u w=0.8u
m18540 2602 2570 VDDREF VDDREF pch l=0.04u w=0.8u
m18541 2603 2571 VDDREF VDDREF pch l=0.04u w=0.8u
m18542 2604 2572 VDDREF VDDREF pch l=0.04u w=0.8u
m18543 2605 2573 VDDREF VDDREF pch l=0.04u w=0.8u
m18544 2606 2574 VDDREF VDDREF pch l=0.04u w=0.8u
m18545 2607 2575 VDDREF VDDREF pch l=0.04u w=0.8u
m18546 2608 2576 VDDREF VDDREF pch l=0.04u w=0.8u
m18547 2609 2577 VDDREF VDDREF pch l=0.04u w=0.8u
m18548 VDDREF 2613 30371 VDDREF pch l=0.04u w=0.12u
m18549 VDDREF 2614 30372 VDDREF pch l=0.04u w=0.12u
m18550 VDDREF 2631 VDDREF VDDREF pch l=0.26u w=1u
m18551 30382 2581 2597 VDDREF pch l=0.04u w=0.12u
m18552 30383 2582 2598 VDDREF pch l=0.04u w=0.12u
m18553 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18554 VDDREF 2641 VDDREF VDDREF pch l=0.26u w=1u
m18555 VDDREF 2642 VDDREF VDDREF pch l=0.26u w=1u
m18556 VDDREF 2645 VDDREF VDDREF pch l=0.26u w=1u
m18557 VDDREF 2646 VDDREF VDDREF pch l=0.26u w=1u
m18558 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18559 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18560 VDDREF 2616 30375 VDDREF pch l=0.04u w=0.12u
m18561 2610 2491 VDDREF VDDREF pch l=0.04u w=0.8u
m18562 2611 2595 VDDREF VDDREF pch l=0.04u w=0.8u
m18563 2496 91 2486 VDDREF pch l=0.04u w=0.8u
m18564 2612 2596 VDDREF VDDREF pch l=0.04u w=0.8u
m18565 2497 2490 2097 VDDREF pch l=0.04u w=0.8u
m18566 2498 2486 FRAC[16] VDDREF pch l=0.04u w=0.8u
m18567 2499 2287 2155 VDDREF pch l=0.04u w=0.8u
m18568 2500 2288 FRAC[16] VDDREF pch l=0.04u w=0.8u
m18569 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18570 2613 2589 VDDREF VDDREF pch l=0.04u w=0.8u
m18571 2614 2590 VDDREF VDDREF pch l=0.04u w=0.8u
m18572 VDDREF 2628 30382 VDDREF pch l=0.04u w=0.12u
m18573 VDDREF 2629 30383 VDDREF pch l=0.04u w=0.12u
m18574 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18575 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18576 2615 5232 VDDREF VDDREF pch l=0.04u w=0.8u
m18577 VDDREF 2652 VDDREF VDDREF pch l=0.26u w=1u
m18578 VDDREF 2655 VDDREF VDDREF pch l=0.26u w=1u
m18579 VDDREF 2656 VDDREF VDDREF pch l=0.26u w=1u
m18580 VDDREF 2659 VDDREF VDDREF pch l=0.26u w=1u
m18581 VDDREF 2660 VDDREF VDDREF pch l=0.26u w=1u
m18582 VDDREF 2663 VDDREF VDDREF pch l=0.26u w=1u
m18583 VDDREF 2664 VDDREF VDDREF pch l=0.26u w=1u
m18584 2616 2593 VDDREF VDDREF pch l=0.04u w=0.8u
m18585 VDDREF 2302 2611 VDDREF pch l=0.04u w=0.8u
m18586 91 2486 2496 VDDREF pch l=0.04u w=0.8u
m18587 VDDREF 2303 2612 VDDREF pch l=0.04u w=0.8u
m18588 2490 2097 2497 VDDREF pch l=0.04u w=0.8u
m18589 2486 FRAC[16] 2498 VDDREF pch l=0.04u w=0.8u
m18590 VDDREF 2631 VDDREF VDDREF pch l=0.26u w=1u
m18591 2287 2155 2499 VDDREF pch l=0.04u w=0.8u
m18592 2288 FRAC[16] 2500 VDDREF pch l=0.04u w=0.8u
m18593 2618 2599 VDDREF VDDREF pch l=0.04u w=0.8u
m18594 2619 2600 VDDREF VDDREF pch l=0.04u w=0.8u
m18595 2620 2602 VDDREF VDDREF pch l=0.04u w=0.8u
m18596 2621 2603 VDDREF VDDREF pch l=0.04u w=0.8u
m18597 2622 2604 VDDREF VDDREF pch l=0.04u w=0.8u
m18598 2623 2605 VDDREF VDDREF pch l=0.04u w=0.8u
m18599 2624 2606 VDDREF VDDREF pch l=0.04u w=0.8u
m18600 2625 2607 VDDREF VDDREF pch l=0.04u w=0.8u
m18601 2626 2608 VDDREF VDDREF pch l=0.04u w=0.8u
m18602 2627 2609 VDDREF VDDREF pch l=0.04u w=0.8u
m18603 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18604 VDDREF 2641 VDDREF VDDREF pch l=0.26u w=1u
m18605 VDDREF 2642 VDDREF VDDREF pch l=0.26u w=1u
m18606 VDDREF 2645 VDDREF VDDREF pch l=0.26u w=1u
m18607 VDDREF 2646 VDDREF VDDREF pch l=0.26u w=1u
m18608 2628 2597 VDDREF VDDREF pch l=0.04u w=0.8u
m18609 2629 2598 VDDREF VDDREF pch l=0.04u w=0.8u
m18610 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18611 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18612 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18613 2617 2630 2491 VDDREF pch l=0.04u w=0.8u
m18614 2611 1370 VDDREF VDDREF pch l=0.04u w=0.8u
m18615 2612 1371 VDDREF VDDREF pch l=0.04u w=0.8u
m18616 2632 2632 VDDREF VDDREF pch l=0.04u w=1u
m18617 VDDREF 2327 2618 VDDREF pch l=0.04u w=0.8u
m18618 VDDREF 2329 2619 VDDREF pch l=0.04u w=0.8u
m18619 VDDREF 2331 2620 VDDREF pch l=0.04u w=0.8u
m18620 VDDREF 2333 2621 VDDREF pch l=0.04u w=0.8u
m18621 VDDREF 2334 2622 VDDREF pch l=0.04u w=0.8u
m18622 VDDREF 2336 2623 VDDREF pch l=0.04u w=0.8u
m18623 VDDREF 2337 2624 VDDREF pch l=0.04u w=0.8u
m18624 VDDREF 2338 2625 VDDREF pch l=0.04u w=0.8u
m18625 VDDREF 2340 2626 VDDREF pch l=0.04u w=0.8u
m18626 VDDREF 2341 2627 VDDREF pch l=0.04u w=0.8u
m18627 2636 2578 2613 VDDREF pch l=0.04u w=0.8u
m18628 2637 2579 2614 VDDREF pch l=0.04u w=0.8u
m18629 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18630 2640 2640 VDDREF VDDREF pch l=0.04u w=1u
m18631 2643 2643 VDDREF VDDREF pch l=0.04u w=1u
m18632 2644 2644 VDDREF VDDREF pch l=0.04u w=1u
m18633 2647 2647 VDDREF VDDREF pch l=0.04u w=1u
m18634 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18635 VDDREF 2652 VDDREF VDDREF pch l=0.26u w=1u
m18636 VDDREF 2655 VDDREF VDDREF pch l=0.26u w=1u
m18637 VDDREF 2656 VDDREF VDDREF pch l=0.26u w=1u
m18638 VDDREF 2659 VDDREF VDDREF pch l=0.26u w=1u
m18639 VDDREF 2660 VDDREF VDDREF pch l=0.26u w=1u
m18640 VDDREF 2663 VDDREF VDDREF pch l=0.26u w=1u
m18641 VDDREF 2664 VDDREF VDDREF pch l=0.26u w=1u
m18642 2648 2759 VDDREF VDDREF pch l=0.04u w=0.8u
m18643 313 2649 VDDREF VDDREF pch l=0.04u w=0.8u
m18644 2630 2491 2617 VDDREF pch l=0.04u w=0.8u
m18645 VDDREF 91 2633 VDDREF pch l=0.04u w=0.8u
m18646 2618 1380 VDDREF VDDREF pch l=0.04u w=0.8u
m18647 VDDREF 2490 2634 VDDREF pch l=0.04u w=0.8u
m18648 2619 1382 VDDREF VDDREF pch l=0.04u w=0.8u
m18649 VDDREF 2486 2635 VDDREF pch l=0.04u w=0.8u
m18650 2620 1384 VDDREF VDDREF pch l=0.04u w=0.8u
m18651 2621 1385 VDDREF VDDREF pch l=0.04u w=0.8u
m18652 2622 1386 VDDREF VDDREF pch l=0.04u w=0.8u
m18653 VDDREF 2287 2638 VDDREF pch l=0.04u w=0.8u
m18654 2623 1387 VDDREF VDDREF pch l=0.04u w=0.8u
m18655 2624 1388 VDDREF VDDREF pch l=0.04u w=0.8u
m18656 2625 1389 VDDREF VDDREF pch l=0.04u w=0.8u
m18657 VDDREF 2288 2639 VDDREF pch l=0.04u w=0.8u
m18658 2626 1390 VDDREF VDDREF pch l=0.04u w=0.8u
m18659 2627 1391 VDDREF VDDREF pch l=0.04u w=0.8u
m18660 30409 4328 2636 VDDREF pch l=0.04u w=0.12u
m18661 30410 4328 2637 VDDREF pch l=0.04u w=0.12u
m18662 VDDREF 2674 VDDREF VDDREF pch l=0.26u w=1u
m18663 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18664 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18665 2650 2581 2628 VDDREF pch l=0.04u w=0.8u
m18666 2651 2582 2629 VDDREF pch l=0.04u w=0.8u
m18667 2653 2653 VDDREF VDDREF pch l=0.04u w=1u
m18668 2654 2654 VDDREF VDDREF pch l=0.04u w=1u
m18669 2657 2657 VDDREF VDDREF pch l=0.04u w=1u
m18670 2658 2658 VDDREF VDDREF pch l=0.04u w=1u
m18671 2661 2661 VDDREF VDDREF pch l=0.04u w=1u
m18672 2662 2662 VDDREF VDDREF pch l=0.04u w=1u
m18673 2665 2665 VDDREF VDDREF pch l=0.04u w=1u
m18674 VDDREF 2759 2648 VDDREF pch l=0.04u w=0.8u
m18675 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18676 30417 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m18677 2667 2525 VDDREF VDDREF pch l=0.04u w=0.8u
m18678 2668 2526 VDDREF VDDREF pch l=0.04u w=0.8u
m18679 VDDREF 2681 30409 VDDREF pch l=0.04u w=0.12u
m18680 VDDREF 2682 30410 VDDREF pch l=0.04u w=0.12u
m18681 2675 2675 VDDREF VDDREF pch l=0.04u w=1u
m18682 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18683 VDDREF 2693 VDDREF VDDREF pch l=0.26u w=1u
m18684 30418 4353 2650 VDDREF pch l=0.04u w=0.12u
m18685 30419 11 2651 VDDREF pch l=0.04u w=0.12u
m18686 2676 2676 VDDREF VDDREF pch l=0.04u w=1u
m18687 2666 2617 30417 VDDREF pch l=0.04u w=0.8u
m18688 2677 2508 VDDREF VDDREF pch l=0.04u w=0.8u
m18689 VDDREF 2611 2667 VDDREF pch l=0.04u w=0.8u
m18690 VDDREF 2612 2668 VDDREF pch l=0.04u w=0.8u
m18691 2669 91 VDDREF VDDREF pch l=0.04u w=0.8u
m18692 2678 2544 VDDREF VDDREF pch l=0.04u w=0.8u
m18693 2670 2490 VDDREF VDDREF pch l=0.04u w=0.8u
m18694 2679 2545 VDDREF VDDREF pch l=0.04u w=0.8u
m18695 2671 2486 VDDREF VDDREF pch l=0.04u w=0.8u
m18696 2680 2546 VDDREF VDDREF pch l=0.04u w=0.8u
m18697 2681 2636 VDDREF VDDREF pch l=0.04u w=0.8u
m18698 2682 2637 VDDREF VDDREF pch l=0.04u w=0.8u
m18699 2683 2547 VDDREF VDDREF pch l=0.04u w=0.8u
m18700 2684 2548 VDDREF VDDREF pch l=0.04u w=0.8u
m18701 2672 2287 VDDREF VDDREF pch l=0.04u w=0.8u
m18702 2685 2549 VDDREF VDDREF pch l=0.04u w=0.8u
m18703 2686 2550 VDDREF VDDREF pch l=0.04u w=0.8u
m18704 2687 2551 VDDREF VDDREF pch l=0.04u w=0.8u
m18705 2673 2288 VDDREF VDDREF pch l=0.04u w=0.8u
m18706 2688 2552 VDDREF VDDREF pch l=0.04u w=0.8u
m18707 2689 2553 VDDREF VDDREF pch l=0.04u w=0.8u
m18708 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18709 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18710 2692 2692 VDDREF VDDREF pch l=0.04u w=1u
m18711 VDDREF 2696 30418 VDDREF pch l=0.04u w=0.12u
m18712 VDDREF 2697 30419 VDDREF pch l=0.04u w=0.12u
m18713 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18714 VDDREF 2197 2677 VDDREF pch l=0.04u w=0.8u
m18715 VDDREF 2486 2669 VDDREF pch l=0.04u w=0.8u
m18716 VDDREF 2618 2678 VDDREF pch l=0.04u w=0.8u
m18717 VDDREF 2704 VDDREF VDDREF pch l=0.26u w=1u
m18718 VDDREF 2097 2670 VDDREF pch l=0.04u w=0.8u
m18719 VDDREF 2619 2679 VDDREF pch l=0.04u w=0.8u
m18720 VDDREF FRAC[16] 2671 VDDREF pch l=0.04u w=0.8u
m18721 VDDREF 2620 2680 VDDREF pch l=0.04u w=0.8u
m18722 VDDREF 2621 2683 VDDREF pch l=0.04u w=0.8u
m18723 VDDREF 2622 2684 VDDREF pch l=0.04u w=0.8u
m18724 VDDREF 2155 2672 VDDREF pch l=0.04u w=0.8u
m18725 VDDREF 2623 2685 VDDREF pch l=0.04u w=0.8u
m18726 VDDREF 2624 2686 VDDREF pch l=0.04u w=0.8u
m18727 VDDREF 2625 2687 VDDREF pch l=0.04u w=0.8u
m18728 VDDREF FRAC[16] 2673 VDDREF pch l=0.04u w=0.8u
m18729 VDDREF 2626 2688 VDDREF pch l=0.04u w=0.8u
m18730 VDDREF 2627 2689 VDDREF pch l=0.04u w=0.8u
m18731 VDDREF 2690 2691 VDDREF pch l=0.04u w=1u
m18732 2696 2650 VDDREF VDDREF pch l=0.04u w=0.8u
m18733 2697 2651 VDDREF VDDREF pch l=0.04u w=0.8u
m18734 2700 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m18735 2701 110 VDDREF VDDREF pch l=0.04u w=0.8u
m18736 293 2702 VDDREF VDDREF pch l=0.04u w=0.8u
m18737 2703 2703 VDDREF VDDREF pch l=0.04u w=1u
m18738 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18739 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18740 2713 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18741 2714 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18742 VDDREF 2695 2694 VDDREF pch l=0.04u w=1u
m18743 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18744 VDDREF 2698 2699 VDDREF pch l=0.04u w=1u
m18745 VDDREF 2197 2700 VDDREF pch l=0.04u w=0.8u
m18746 2717 2197 VDDREF VDDREF pch l=0.04u w=0.8u
m18747 VDDREF 125 2701 VDDREF pch l=0.04u w=0.8u
m18748 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m18749 VDDREF 2705 2706 VDDREF pch l=0.04u w=1u
m18750 VDDREF 2708 2707 VDDREF pch l=0.04u w=1u
m18751 2466 2753 VDDREF VDDREF pch l=0.04u w=0.8u
m18752 2718 2795 VDDREF VDDREF pch l=0.04u w=0.8u
m18753 2468 2754 VDDREF VDDREF pch l=0.04u w=0.8u
m18754 2723 1853 VDDREF VDDREF pch l=0.04u w=0.8u
m18755 2724 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m18756 2725 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m18757 VDDREF 2709 2710 VDDREF pch l=0.04u w=1u
m18758 VDDREF 2712 2711 VDDREF pch l=0.04u w=1u
m18759 2470 2755 VDDREF VDDREF pch l=0.04u w=0.8u
m18760 2726 FRAC[8] VDDREF VDDREF pch l=0.04u w=0.8u
m18761 VDDREF 2774 2715 VDDREF pch l=0.04u w=0.8u
m18762 2727 2796 VDDREF VDDREF pch l=0.04u w=0.8u
m18763 2728 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18764 2729 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18765 2730 2804 VDDREF VDDREF pch l=0.04u w=0.8u
m18766 2474 2757 VDDREF VDDREF pch l=0.04u w=0.8u
m18767 2731 2805 VDDREF VDDREF pch l=0.04u w=0.8u
m18768 2732 2715 VDDREF VDDREF pch l=0.04u w=0.8u
m18769 2733 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18770 2734 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18771 2735 2808 VDDREF VDDREF pch l=0.04u w=0.8u
m18772 2478 2758 VDDREF VDDREF pch l=0.04u w=0.8u
m18773 2736 FRAC[8] VDDREF VDDREF pch l=0.04u w=0.8u
m18774 2737 2715 VDDREF VDDREF pch l=0.04u w=0.8u
m18775 2738 PD VDDREF VDDREF pch l=0.04u w=0.8u
m18776 VDDREF 2746 2716 VDDREF pch l=0.04u w=0.8u
m18777 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18778 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18779 VDDREF 2889 2466 VDDREF pch l=0.04u w=0.8u
m18780 VDDREF 2793 2718 VDDREF pch l=0.04u w=0.8u
m18781 VDDREF 2719 2720 VDDREF pch l=0.04u w=1u
m18782 VDDREF 2722 2721 VDDREF pch l=0.04u w=1u
m18783 VDDREF 2890 2468 VDDREF pch l=0.04u w=0.8u
m18784 VDDREF 2794 2723 VDDREF pch l=0.04u w=0.8u
m18785 VDDREF 2928 2724 VDDREF pch l=0.04u w=0.8u
m18786 VDDREF 2929 2725 VDDREF pch l=0.04u w=0.8u
m18787 VDDREF 2891 2470 VDDREF pch l=0.04u w=0.8u
m18788 VDDREF 2795 2726 VDDREF pch l=0.04u w=0.8u
m18789 VDDREF 131 2727 VDDREF pch l=0.04u w=0.8u
m18790 VDDREF 2796 2730 VDDREF pch l=0.04u w=0.8u
m18791 VDDREF 2892 2474 VDDREF pch l=0.04u w=0.8u
m18792 VDDREF 2797 2731 VDDREF pch l=0.04u w=0.8u
m18793 VDDREF 2798 2732 VDDREF pch l=0.04u w=0.8u
m18794 VDDREF 2799 2735 VDDREF pch l=0.04u w=0.8u
m18795 VDDREF 2893 2478 VDDREF pch l=0.04u w=0.8u
m18796 VDDREF 2800 2736 VDDREF pch l=0.04u w=0.8u
m18797 VDDREF FBDIV[8] 2737 VDDREF pch l=0.04u w=0.8u
m18798 2740 4328 2681 VDDREF pch l=0.04u w=0.8u
m18799 2741 4328 2682 VDDREF pch l=0.04u w=0.8u
m18800 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m18801 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18802 VDDREF 2858 VDDREF VDDREF pch l=0.26u w=1u
m18803 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m18804 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m18805 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m18806 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m18807 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m18808 2747 2700 VDDREF VDDREF pch l=0.04u w=0.8u
m18809 2739 2508 2197 VDDREF pch l=0.04u w=0.8u
m18810 2748 125 VDDREF VDDREF pch l=0.04u w=0.8u
m18811 30481 2713 2740 VDDREF pch l=0.04u w=0.12u
m18812 30482 2714 2741 VDDREF pch l=0.04u w=0.12u
m18813 2756 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18814 2749 4328 2742 VDDREF pch l=0.04u w=0.8u
m18815 2750 4328 2743 VDDREF pch l=0.04u w=0.8u
m18816 2751 4328 2744 VDDREF pch l=0.04u w=0.8u
m18817 2752 4328 2745 VDDREF pch l=0.04u w=0.8u
m18818 2759 2738 VDDREF VDDREF pch l=0.04u w=0.8u
m18819 VDDREF 5232 2746 VDDREF pch l=0.04u w=0.4u
m18820 VDDREF 2775 VDDREF VDDREF pch l=0.26u w=1u
m18821 VDDREF 2778 VDDREF VDDREF pch l=0.26u w=1u
m18822 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m18823 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m18824 2508 2197 2739 VDDREF pch l=0.04u w=0.8u
m18825 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m18826 VDDREF 3737 2753 VDDREF pch l=0.04u w=0.8u
m18827 2762 2793 VDDREF VDDREF pch l=0.04u w=0.8u
m18828 VDDREF 3739 2754 VDDREF pch l=0.04u w=0.8u
m18829 2763 2794 VDDREF VDDREF pch l=0.04u w=0.8u
m18830 2764 2724 VDDREF VDDREF pch l=0.04u w=0.8u
m18831 2765 2725 VDDREF VDDREF pch l=0.04u w=0.8u
m18832 VDDREF 3741 2755 VDDREF pch l=0.04u w=0.8u
m18833 2766 2795 VDDREF VDDREF pch l=0.04u w=0.8u
m18834 VDDREF 2783 30481 VDDREF pch l=0.04u w=0.12u
m18835 VDDREF 2784 30482 VDDREF pch l=0.04u w=0.12u
m18836 2767 131 VDDREF VDDREF pch l=0.04u w=0.8u
m18837 30490 2728 2749 VDDREF pch l=0.04u w=0.12u
m18838 30491 2729 2750 VDDREF pch l=0.04u w=0.12u
m18839 2768 2796 VDDREF VDDREF pch l=0.04u w=0.8u
m18840 VDDREF 3745 2757 VDDREF pch l=0.04u w=0.8u
m18841 2769 2797 VDDREF VDDREF pch l=0.04u w=0.8u
m18842 2770 2798 VDDREF VDDREF pch l=0.04u w=0.8u
m18843 30492 2733 2751 VDDREF pch l=0.04u w=0.12u
m18844 30493 2734 2752 VDDREF pch l=0.04u w=0.12u
m18845 2771 2799 VDDREF VDDREF pch l=0.04u w=0.8u
m18846 VDDREF 3749 2758 VDDREF pch l=0.04u w=0.8u
m18847 2772 2800 VDDREF VDDREF pch l=0.04u w=0.8u
m18848 2773 FBDIV[8] VDDREF VDDREF pch l=0.04u w=0.8u
m18849 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18850 VDDREF 2696 2759 VDDREF pch l=0.04u w=0.8u
m18851 2746 5232 VDDREF VDDREF pch l=0.04u w=0.4u
m18852 VDDREF 2858 VDDREF VDDREF pch l=0.26u w=1u
m18853 2776 2776 VDDREF VDDREF pch l=0.04u w=1u
m18854 2777 2777 VDDREF VDDREF pch l=0.04u w=1u
m18855 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m18856 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m18857 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m18858 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m18859 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m18860 2761 110 125 VDDREF pch l=0.04u w=0.8u
m18861 2753 2947 VDDREF VDDREF pch l=0.04u w=0.8u
m18862 2754 2948 VDDREF VDDREF pch l=0.04u w=0.8u
m18863 2755 2949 VDDREF VDDREF pch l=0.04u w=0.8u
m18864 2783 2740 VDDREF VDDREF pch l=0.04u w=0.8u
m18865 2784 2741 VDDREF VDDREF pch l=0.04u w=0.8u
m18866 VDDREF 2802 30490 VDDREF pch l=0.04u w=0.12u
m18867 VDDREF 2803 30491 VDDREF pch l=0.04u w=0.12u
m18868 2757 2950 VDDREF VDDREF pch l=0.04u w=0.8u
m18869 VDDREF 2806 30492 VDDREF pch l=0.04u w=0.12u
m18870 VDDREF 2807 30493 VDDREF pch l=0.04u w=0.12u
m18871 2758 2951 VDDREF VDDREF pch l=0.04u w=0.8u
m18872 2785 4328 2774 VDDREF pch l=0.04u w=0.8u
m18873 2759 2697 VDDREF VDDREF pch l=0.04u w=0.8u
m18874 VDDREF 2738 2746 VDDREF pch l=0.04u w=0.12u
m18875 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m18876 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m18877 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m18878 2779 2739 VDDREF VDDREF pch l=0.04u w=0.8u
m18879 110 125 2761 VDDREF pch l=0.04u w=0.8u
m18880 VDDREF 2816 2753 VDDREF pch l=0.04u w=0.8u
m18881 VDDREF 2817 2754 VDDREF pch l=0.04u w=0.8u
m18882 VDDREF 2818 2755 VDDREF pch l=0.04u w=0.8u
m18883 2802 2749 VDDREF VDDREF pch l=0.04u w=0.8u
m18884 2803 2750 VDDREF VDDREF pch l=0.04u w=0.8u
m18885 VDDREF 2819 2757 VDDREF pch l=0.04u w=0.8u
m18886 2806 2751 VDDREF VDDREF pch l=0.04u w=0.8u
m18887 2807 2752 VDDREF VDDREF pch l=0.04u w=0.8u
m18888 VDDREF 2820 2758 VDDREF pch l=0.04u w=0.8u
m18889 2809 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18890 2810 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18891 2780 2795 2793 VDDREF pch l=0.04u w=0.8u
m18892 2781 1853 2794 VDDREF pch l=0.04u w=0.8u
m18893 2811 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18894 2812 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m18895 2782 FRAC[8] 2795 VDDREF pch l=0.04u w=0.8u
m18896 30505 2756 2785 VDDREF pch l=0.04u w=0.12u
m18897 2786 2796 131 VDDREF pch l=0.04u w=0.8u
m18898 2787 2804 2796 VDDREF pch l=0.04u w=0.8u
m18899 2788 2805 2797 VDDREF pch l=0.04u w=0.8u
m18900 2789 2715 2798 VDDREF pch l=0.04u w=0.8u
m18901 2790 2808 2799 VDDREF pch l=0.04u w=0.8u
m18902 2791 FRAC[8] 2800 VDDREF pch l=0.04u w=0.8u
m18903 2792 2715 FBDIV[8] VDDREF pch l=0.04u w=0.8u
m18904 VDDREF 2822 VDDREF VDDREF pch l=0.26u w=1u
m18905 VDDREF 2858 VDDREF VDDREF pch l=0.26u w=1u
m18906 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m18907 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m18908 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m18909 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m18910 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m18911 VDDREF 2583 2779 VDDREF pch l=0.04u w=0.8u
m18912 2795 2793 2780 VDDREF pch l=0.04u w=0.8u
m18913 1853 2794 2781 VDDREF pch l=0.04u w=0.8u
m18914 FRAC[8] 2795 2782 VDDREF pch l=0.04u w=0.8u
m18915 2813 2713 2783 VDDREF pch l=0.04u w=0.8u
m18916 2814 2714 2784 VDDREF pch l=0.04u w=0.8u
m18917 VDDREF 2833 30505 VDDREF pch l=0.04u w=0.12u
m18918 2796 131 2786 VDDREF pch l=0.04u w=0.8u
m18919 2804 2796 2787 VDDREF pch l=0.04u w=0.8u
m18920 2805 2797 2788 VDDREF pch l=0.04u w=0.8u
m18921 2715 2798 2789 VDDREF pch l=0.04u w=0.8u
m18922 2808 2799 2790 VDDREF pch l=0.04u w=0.8u
m18923 FRAC[8] 2800 2791 VDDREF pch l=0.04u w=0.8u
m18924 2715 FBDIV[8] 2792 VDDREF pch l=0.04u w=0.8u
m18925 2821 2821 VDDREF VDDREF pch l=0.04u w=1u
m18926 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m18927 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m18928 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m18929 2815 2761 VDDREF VDDREF pch l=0.04u w=0.8u
m18930 VDDREF 2845 2816 VDDREF pch l=0.04u w=0.8u
m18931 VDDREF 2846 2817 VDDREF pch l=0.04u w=0.8u
m18932 VDDREF 2847 2818 VDDREF pch l=0.04u w=0.8u
m18933 30526 4328 2813 VDDREF pch l=0.04u w=0.12u
m18934 30527 4328 2814 VDDREF pch l=0.04u w=0.12u
m18935 2833 2785 VDDREF VDDREF pch l=0.04u w=0.8u
m18936 2825 2728 2802 VDDREF pch l=0.04u w=0.8u
m18937 2826 2729 2803 VDDREF pch l=0.04u w=0.8u
m18938 VDDREF 2848 2819 VDDREF pch l=0.04u w=0.8u
m18939 2827 2733 2806 VDDREF pch l=0.04u w=0.8u
m18940 2828 2734 2807 VDDREF pch l=0.04u w=0.8u
m18941 VDDREF 2849 2820 VDDREF pch l=0.04u w=0.8u
m18942 2829 4328 2823 VDDREF pch l=0.04u w=0.8u
m18943 2830 4328 2824 VDDREF pch l=0.04u w=0.8u
m18944 2831 4328 2764 VDDREF pch l=0.04u w=0.8u
m18945 2832 4328 2765 VDDREF pch l=0.04u w=0.8u
m18946 VDDREF 2858 VDDREF VDDREF pch l=0.26u w=1u
m18947 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m18948 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m18949 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m18950 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m18951 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m18952 2844 2779 VDDREF VDDREF pch l=0.04u w=0.8u
m18953 VDDREF 2667 2815 VDDREF pch l=0.04u w=0.8u
m18954 VDDREF 2851 30526 VDDREF pch l=0.04u w=0.12u
m18955 VDDREF 2852 30527 VDDREF pch l=0.04u w=0.12u
m18956 30545 4328 2825 VDDREF pch l=0.04u w=0.12u
m18957 30546 4328 2826 VDDREF pch l=0.04u w=0.12u
m18958 30547 4328 2827 VDDREF pch l=0.04u w=0.12u
m18959 30548 4328 2828 VDDREF pch l=0.04u w=0.12u
m18960 30551 2809 2829 VDDREF pch l=0.04u w=0.12u
m18961 30552 2810 2830 VDDREF pch l=0.04u w=0.12u
m18962 2834 2780 VDDREF VDDREF pch l=0.04u w=0.8u
m18963 2835 2781 VDDREF VDDREF pch l=0.04u w=0.8u
m18964 30553 2811 2831 VDDREF pch l=0.04u w=0.12u
m18965 30554 2812 2832 VDDREF pch l=0.04u w=0.12u
m18966 2836 2782 VDDREF VDDREF pch l=0.04u w=0.8u
m18967 2837 2786 VDDREF VDDREF pch l=0.04u w=0.8u
m18968 2838 2787 VDDREF VDDREF pch l=0.04u w=0.8u
m18969 2839 2788 VDDREF VDDREF pch l=0.04u w=0.8u
m18970 2840 2789 VDDREF VDDREF pch l=0.04u w=0.8u
m18971 2841 2790 VDDREF VDDREF pch l=0.04u w=0.8u
m18972 2842 2791 VDDREF VDDREF pch l=0.04u w=0.8u
m18973 2843 2792 VDDREF VDDREF pch l=0.04u w=0.8u
m18974 2850 155 VDDREF VDDREF pch l=0.04u w=0.8u
m18975 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m18976 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m18977 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m18978 VDDREF 2677 2844 VDDREF pch l=0.04u w=0.8u
m18979 2851 2813 VDDREF VDDREF pch l=0.04u w=0.8u
m18980 2852 2814 VDDREF VDDREF pch l=0.04u w=0.8u
m18981 VDDREF 2854 30545 VDDREF pch l=0.04u w=0.12u
m18982 VDDREF 2855 30546 VDDREF pch l=0.04u w=0.12u
m18983 VDDREF 2856 30547 VDDREF pch l=0.04u w=0.12u
m18984 VDDREF 2857 30548 VDDREF pch l=0.04u w=0.12u
m18985 VDDREF 2858 VDDREF VDDREF pch l=0.26u w=1u
m18986 VDDREF 2861 30551 VDDREF pch l=0.04u w=0.12u
m18987 VDDREF 2862 30552 VDDREF pch l=0.04u w=0.12u
m18988 VDDREF 3228 2845 VDDREF pch l=0.04u w=0.8u
m18989 VDDREF 2678 2834 VDDREF pch l=0.04u w=0.8u
m18990 VDDREF 3229 2846 VDDREF pch l=0.04u w=0.8u
m18991 VDDREF 2679 2835 VDDREF pch l=0.04u w=0.8u
m18992 VDDREF 2863 30553 VDDREF pch l=0.04u w=0.12u
m18993 VDDREF 2864 30554 VDDREF pch l=0.04u w=0.12u
m18994 VDDREF 3230 2847 VDDREF pch l=0.04u w=0.8u
m18995 VDDREF 2680 2836 VDDREF pch l=0.04u w=0.8u
m18996 2853 2756 2833 VDDREF pch l=0.04u w=0.8u
m18997 VDDREF 2683 2837 VDDREF pch l=0.04u w=0.8u
m18998 VDDREF 2684 2838 VDDREF pch l=0.04u w=0.8u
m18999 VDDREF 3231 2848 VDDREF pch l=0.04u w=0.8u
m19000 VDDREF 2685 2839 VDDREF pch l=0.04u w=0.8u
m19001 VDDREF 2686 2840 VDDREF pch l=0.04u w=0.8u
m19002 VDDREF 2687 2841 VDDREF pch l=0.04u w=0.8u
m19003 VDDREF 3232 2849 VDDREF pch l=0.04u w=0.8u
m19004 VDDREF 2688 2842 VDDREF pch l=0.04u w=0.8u
m19005 VDDREF 2689 2843 VDDREF pch l=0.04u w=0.8u
m19006 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m19007 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m19008 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m19009 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m19010 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m19011 2854 2825 VDDREF VDDREF pch l=0.04u w=0.8u
m19012 2855 2826 VDDREF VDDREF pch l=0.04u w=0.8u
m19013 2856 2827 VDDREF VDDREF pch l=0.04u w=0.8u
m19014 2857 2828 VDDREF VDDREF pch l=0.04u w=0.8u
m19015 2859 2859 VDDREF VDDREF pch l=0.04u w=1u
m19016 2860 2815 VDDREF VDDREF pch l=0.04u w=0.8u
m19017 2861 2829 VDDREF VDDREF pch l=0.04u w=0.8u
m19018 2862 2830 VDDREF VDDREF pch l=0.04u w=0.8u
m19019 2845 3500 VDDREF VDDREF pch l=0.04u w=0.8u
m19020 2846 3501 VDDREF VDDREF pch l=0.04u w=0.8u
m19021 2863 2831 VDDREF VDDREF pch l=0.04u w=0.8u
m19022 2864 2832 VDDREF VDDREF pch l=0.04u w=0.8u
m19023 2847 3502 VDDREF VDDREF pch l=0.04u w=0.8u
m19024 30579 4328 2853 VDDREF pch l=0.04u w=0.12u
m19025 2848 3503 VDDREF VDDREF pch l=0.04u w=0.8u
m19026 2849 3504 VDDREF VDDREF pch l=0.04u w=0.8u
m19027 2865 155 VDDREF VDDREF pch l=0.04u w=0.8u
m19028 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m19029 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m19030 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m19031 2866 2739 VDDREF VDDREF pch l=0.04u w=0.8u
m19032 VDDREF 2701 2860 VDDREF pch l=0.04u w=0.8u
m19033 VDDREF 3777 2845 VDDREF pch l=0.04u w=0.8u
m19034 VDDREF 3778 2846 VDDREF pch l=0.04u w=0.8u
m19035 VDDREF 3779 2847 VDDREF pch l=0.04u w=0.8u
m19036 2867 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19037 2868 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19038 VDDREF 2884 30579 VDDREF pch l=0.04u w=0.12u
m19039 VDDREF 3780 2848 VDDREF pch l=0.04u w=0.8u
m19040 VDDREF 3781 2849 VDDREF pch l=0.04u w=0.8u
m19041 2869 2834 VDDREF VDDREF pch l=0.04u w=0.8u
m19042 2870 2835 VDDREF VDDREF pch l=0.04u w=0.8u
m19043 2871 2836 VDDREF VDDREF pch l=0.04u w=0.8u
m19044 2872 2837 VDDREF VDDREF pch l=0.04u w=0.8u
m19045 2873 2838 VDDREF VDDREF pch l=0.04u w=0.8u
m19046 2874 2839 VDDREF VDDREF pch l=0.04u w=0.8u
m19047 2875 2840 VDDREF VDDREF pch l=0.04u w=0.8u
m19048 2876 2841 VDDREF VDDREF pch l=0.04u w=0.8u
m19049 2877 2842 VDDREF VDDREF pch l=0.04u w=0.8u
m19050 2878 2843 VDDREF VDDREF pch l=0.04u w=0.8u
m19051 VDDREF FBDIV[8] 2865 VDDREF pch l=0.04u w=0.8u
m19052 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m19053 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m19054 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m19055 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m19056 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m19057 2884 2853 VDDREF VDDREF pch l=0.04u w=0.8u
m19058 2885 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19059 2886 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19060 2887 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19061 2888 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19062 2880 2809 2861 VDDREF pch l=0.04u w=0.8u
m19063 2881 2810 2862 VDDREF pch l=0.04u w=0.8u
m19064 VDDREF 2718 2869 VDDREF pch l=0.04u w=0.8u
m19065 VDDREF 2723 2870 VDDREF pch l=0.04u w=0.8u
m19066 2882 2811 2863 VDDREF pch l=0.04u w=0.8u
m19067 2883 2812 2864 VDDREF pch l=0.04u w=0.8u
m19068 VDDREF 2726 2871 VDDREF pch l=0.04u w=0.8u
m19069 VDDREF 2727 2872 VDDREF pch l=0.04u w=0.8u
m19070 VDDREF 2730 2873 VDDREF pch l=0.04u w=0.8u
m19071 VDDREF 2731 2874 VDDREF pch l=0.04u w=0.8u
m19072 VDDREF 2732 2875 VDDREF pch l=0.04u w=0.8u
m19073 VDDREF 2735 2876 VDDREF pch l=0.04u w=0.8u
m19074 VDDREF 2736 2877 VDDREF pch l=0.04u w=0.8u
m19075 VDDREF 2737 2878 VDDREF pch l=0.04u w=0.8u
m19076 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m19077 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m19078 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m19079 2896 2926 VDDREF VDDREF pch l=0.04u w=0.8u
m19080 2879 2583 2739 VDDREF pch l=0.04u w=0.8u
m19081 2897 2761 VDDREF VDDREF pch l=0.04u w=0.8u
m19082 30623 4328 2880 VDDREF pch l=0.04u w=0.12u
m19083 30624 4328 2881 VDDREF pch l=0.04u w=0.12u
m19084 VDDREF 2995 2889 VDDREF pch l=0.04u w=0.8u
m19085 VDDREF 2997 2890 VDDREF pch l=0.04u w=0.8u
m19086 30625 4328 2882 VDDREF pch l=0.04u w=0.12u
m19087 30626 4328 2883 VDDREF pch l=0.04u w=0.12u
m19088 VDDREF 3001 2891 VDDREF pch l=0.04u w=0.8u
m19089 2894 4328 2851 VDDREF pch l=0.04u w=0.8u
m19090 2895 4328 2852 VDDREF pch l=0.04u w=0.8u
m19091 VDDREF 3005 2892 VDDREF pch l=0.04u w=0.8u
m19092 VDDREF 3009 2893 VDDREF pch l=0.04u w=0.8u
m19093 VDDREF 2907 VDDREF VDDREF pch l=0.26u w=1u
m19094 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m19095 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m19096 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m19097 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m19098 2901 2850 VDDREF VDDREF pch l=0.04u w=0.8u
m19099 VDDREF 2926 2896 VDDREF pch l=0.04u w=0.8u
m19100 2583 2739 2879 VDDREF pch l=0.04u w=0.8u
m19101 VDDREF 2924 30623 VDDREF pch l=0.04u w=0.12u
m19102 VDDREF 2793 30624 VDDREF pch l=0.04u w=0.12u
m19103 VDDREF 2925 30625 VDDREF pch l=0.04u w=0.12u
m19104 VDDREF 2795 30626 VDDREF pch l=0.04u w=0.12u
m19105 30640 2867 2894 VDDREF pch l=0.04u w=0.12u
m19106 30641 2868 2895 VDDREF pch l=0.04u w=0.12u
m19107 2902 4328 2898 VDDREF pch l=0.04u w=0.8u
m19108 2903 4328 2899 VDDREF pch l=0.04u w=0.8u
m19109 2904 4328 2900 VDDREF pch l=0.04u w=0.8u
m19110 2905 4328 2798 VDDREF pch l=0.04u w=0.8u
m19111 2908 2908 VDDREF VDDREF pch l=0.04u w=1u
m19112 2910 2780 VDDREF VDDREF pch l=0.04u w=0.8u
m19113 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m19114 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m19115 2912 2781 VDDREF VDDREF pch l=0.04u w=0.8u
m19116 2914 2782 VDDREF VDDREF pch l=0.04u w=0.8u
m19117 2915 2786 VDDREF VDDREF pch l=0.04u w=0.8u
m19118 2916 2787 VDDREF VDDREF pch l=0.04u w=0.8u
m19119 2918 2788 VDDREF VDDREF pch l=0.04u w=0.8u
m19120 2919 2789 VDDREF VDDREF pch l=0.04u w=0.8u
m19121 2920 2790 VDDREF VDDREF pch l=0.04u w=0.8u
m19122 2922 2791 VDDREF VDDREF pch l=0.04u w=0.8u
m19123 2923 2792 VDDREF VDDREF pch l=0.04u w=0.8u
m19124 VDDREF 2884 2901 VDDREF pch l=0.04u w=0.8u
m19125 VDDREF 2935 VDDREF VDDREF pch l=0.26u w=1u
m19126 2924 2880 VDDREF VDDREF pch l=0.04u w=0.8u
m19127 2793 2881 VDDREF VDDREF pch l=0.04u w=0.8u
m19128 VDDREF 2936 VDDREF VDDREF pch l=0.26u w=1u
m19129 VDDREF 2939 VDDREF VDDREF pch l=0.26u w=1u
m19130 2925 2882 VDDREF VDDREF pch l=0.04u w=0.8u
m19131 2795 2883 VDDREF VDDREF pch l=0.04u w=0.8u
m19132 VDDREF 2940 VDDREF VDDREF pch l=0.26u w=1u
m19133 VDDREF 2943 VDDREF VDDREF pch l=0.26u w=1u
m19134 VDDREF 2944 30640 VDDREF pch l=0.04u w=0.12u
m19135 VDDREF 2945 30641 VDDREF pch l=0.04u w=0.12u
m19136 30687 2885 2902 VDDREF pch l=0.04u w=0.12u
m19137 30688 2886 2903 VDDREF pch l=0.04u w=0.12u
m19138 30689 2887 2904 VDDREF pch l=0.04u w=0.12u
m19139 30690 2888 2905 VDDREF pch l=0.04u w=0.12u
m19140 30691 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m19141 2906 2667 2761 VDDREF pch l=0.04u w=0.8u
m19142 2823 2947 2909 VDDREF pch l=0.04u w=0.8u
m19143 2928 2948 2911 VDDREF pch l=0.04u w=0.8u
m19144 2930 2949 2913 VDDREF pch l=0.04u w=0.8u
m19145 2743 2950 2917 VDDREF pch l=0.04u w=0.8u
m19146 2745 2951 2921 VDDREF pch l=0.04u w=0.8u
m19147 2934 2934 VDDREF VDDREF pch l=0.04u w=1u
m19148 2937 2937 VDDREF VDDREF pch l=0.04u w=1u
m19149 2938 2938 VDDREF VDDREF pch l=0.04u w=1u
m19150 VDDREF 2956 VDDREF VDDREF pch l=0.26u w=1u
m19151 VDDREF 2959 VDDREF VDDREF pch l=0.26u w=1u
m19152 2941 2941 VDDREF VDDREF pch l=0.04u w=1u
m19153 2942 2942 VDDREF VDDREF pch l=0.04u w=1u
m19154 2944 2894 VDDREF VDDREF pch l=0.04u w=0.8u
m19155 2945 2895 VDDREF VDDREF pch l=0.04u w=0.8u
m19156 VDDREF 2960 30687 VDDREF pch l=0.04u w=0.12u
m19157 VDDREF 2961 30688 VDDREF pch l=0.04u w=0.12u
m19158 VDDREF 2962 30689 VDDREF pch l=0.04u w=0.12u
m19159 VDDREF 2963 30690 VDDREF pch l=0.04u w=0.12u
m19160 VDDREF 2977 2926 VDDREF pch l=0.04u w=0.8u
m19161 2927 2879 30691 VDDREF pch l=0.04u w=0.8u
m19162 2946 2508 VDDREF VDDREF pch l=0.04u w=0.8u
m19163 2667 2761 2906 VDDREF pch l=0.04u w=0.8u
m19164 2947 2909 2823 VDDREF pch l=0.04u w=0.8u
m19165 2948 2911 2928 VDDREF pch l=0.04u w=0.8u
m19166 2949 2913 2930 VDDREF pch l=0.04u w=0.8u
m19167 2950 2917 2743 VDDREF pch l=0.04u w=0.8u
m19168 2951 2921 2745 VDDREF pch l=0.04u w=0.8u
m19169 VDDREF 2932 2933 VDDREF pch l=0.04u w=1u
m19170 2824 2678 2780 VDDREF pch l=0.04u w=0.8u
m19171 2929 2679 2781 VDDREF pch l=0.04u w=0.8u
m19172 2794 2680 2782 VDDREF pch l=0.04u w=0.8u
m19173 2774 2683 2786 VDDREF pch l=0.04u w=0.8u
m19174 2899 2684 2787 VDDREF pch l=0.04u w=0.8u
m19175 2931 2685 2788 VDDREF pch l=0.04u w=0.8u
m19176 2804 2686 2789 VDDREF pch l=0.04u w=0.8u
m19177 2798 2687 2790 VDDREF pch l=0.04u w=0.8u
m19178 2805 2688 2791 VDDREF pch l=0.04u w=0.8u
m19179 2808 2689 2792 VDDREF pch l=0.04u w=0.8u
m19180 2952 2901 VDDREF VDDREF pch l=0.04u w=0.8u
m19181 2955 2896 VDDREF VDDREF pch l=0.04u w=0.8u
m19182 2957 2957 VDDREF VDDREF pch l=0.04u w=1u
m19183 2958 2958 VDDREF VDDREF pch l=0.04u w=1u
m19184 2960 2902 VDDREF VDDREF pch l=0.04u w=0.8u
m19185 2961 2903 VDDREF VDDREF pch l=0.04u w=0.8u
m19186 2962 2904 VDDREF VDDREF pch l=0.04u w=0.8u
m19187 2963 2905 VDDREF VDDREF pch l=0.04u w=0.8u
m19188 30711 2926 VDDREF VDDREF pch l=0.04u w=0.12u
m19189 VDDREF 2465 2946 VDDREF pch l=0.04u w=0.8u
m19190 2678 2780 2824 VDDREF pch l=0.04u w=0.8u
m19191 2679 2781 2929 VDDREF pch l=0.04u w=0.8u
m19192 2680 2782 2794 VDDREF pch l=0.04u w=0.8u
m19193 2683 2786 2774 VDDREF pch l=0.04u w=0.8u
m19194 2684 2787 2899 VDDREF pch l=0.04u w=0.8u
m19195 2685 2788 2931 VDDREF pch l=0.04u w=0.8u
m19196 2686 2789 2804 VDDREF pch l=0.04u w=0.8u
m19197 2687 2790 2798 VDDREF pch l=0.04u w=0.8u
m19198 2688 2791 2805 VDDREF pch l=0.04u w=0.8u
m19199 2689 2792 2808 VDDREF pch l=0.04u w=0.8u
m19200 VDDREF 2865 2952 VDDREF pch l=0.04u w=0.8u
m19201 VDDREF 2954 2953 VDDREF pch l=0.04u w=1u
m19202 VDDREF 3565 2955 VDDREF pch l=0.04u w=0.8u
m19203 2969 3013 VDDREF VDDREF pch l=0.04u w=0.8u
m19204 2970 2969 VDDREF VDDREF pch l=0.04u w=0.8u
m19205 2977 4251 30711 VDDREF pch l=0.04u w=0.12u
m19206 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19207 2971 2867 2944 VDDREF pch l=0.04u w=0.8u
m19208 2972 2868 2945 VDDREF pch l=0.04u w=0.8u
m19209 2978 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m19210 2979 110 VDDREF VDDREF pch l=0.04u w=0.8u
m19211 VDDREF 2947 2964 VDDREF pch l=0.04u w=0.8u
m19212 VDDREF 2948 2965 VDDREF pch l=0.04u w=0.8u
m19213 VDDREF 2949 2966 VDDREF pch l=0.04u w=0.8u
m19214 VDDREF 2950 2967 VDDREF pch l=0.04u w=0.8u
m19215 VDDREF 2951 2968 VDDREF pch l=0.04u w=0.8u
m19216 2955 4064 VDDREF VDDREF pch l=0.04u w=0.8u
m19217 VDDREF 3013 2969 VDDREF pch l=0.04u w=0.8u
m19218 VDDREF 3484 2970 VDDREF pch l=0.04u w=0.8u
m19219 2993 3085 2977 VDDREF pch l=0.04u w=0.8u
m19220 VDDREF 2973 2974 VDDREF pch l=0.04u w=1u
m19221 VDDREF 2976 2975 VDDREF pch l=0.04u w=1u
m19222 30736 4328 2971 VDDREF pch l=0.04u w=0.12u
m19223 30737 4328 2972 VDDREF pch l=0.04u w=0.12u
m19224 2989 2885 2960 VDDREF pch l=0.04u w=0.8u
m19225 2990 2886 2961 VDDREF pch l=0.04u w=0.8u
m19226 2991 2887 2962 VDDREF pch l=0.04u w=0.8u
m19227 2992 2888 2963 VDDREF pch l=0.04u w=0.8u
m19228 VDDREF 2465 2978 VDDREF pch l=0.04u w=0.8u
m19229 2994 2465 VDDREF VDDREF pch l=0.04u w=0.8u
m19230 VDDREF 437 2979 VDDREF pch l=0.04u w=0.8u
m19231 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19232 VDDREF 2980 2981 VDDREF pch l=0.04u w=1u
m19233 VDDREF 2983 2982 VDDREF pch l=0.04u w=1u
m19234 2996 3065 VDDREF VDDREF pch l=0.04u w=0.8u
m19235 2998 1877 VDDREF VDDREF pch l=0.04u w=0.8u
m19236 2999 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m19237 3000 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m19238 VDDREF 2984 2985 VDDREF pch l=0.04u w=1u
m19239 VDDREF 2987 2986 VDDREF pch l=0.04u w=1u
m19240 3002 FRAC[9] VDDREF VDDREF pch l=0.04u w=0.8u
m19241 VDDREF 3038 2988 VDDREF pch l=0.04u w=0.8u
m19242 3003 3066 VDDREF VDDREF pch l=0.04u w=0.8u
m19243 3004 3078 VDDREF VDDREF pch l=0.04u w=0.8u
m19244 3006 2900 VDDREF VDDREF pch l=0.04u w=0.8u
m19245 3007 2988 VDDREF VDDREF pch l=0.04u w=0.8u
m19246 3008 3079 VDDREF VDDREF pch l=0.04u w=0.8u
m19247 3010 FRAC[9] VDDREF VDDREF pch l=0.04u w=0.8u
m19248 3011 2988 VDDREF VDDREF pch l=0.04u w=0.8u
m19249 3012 3062 VDDREF VDDREF pch l=0.04u w=0.8u
m19250 2970 3953 VDDREF VDDREF pch l=0.04u w=0.8u
m19251 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19252 VDDREF 1146 30736 VDDREF pch l=0.04u w=0.12u
m19253 VDDREF 3018 30737 VDDREF pch l=0.04u w=0.12u
m19254 30747 4328 2989 VDDREF pch l=0.04u w=0.12u
m19255 30748 4328 2990 VDDREF pch l=0.04u w=0.12u
m19256 30749 4328 2991 VDDREF pch l=0.04u w=0.12u
m19257 30750 4328 2992 VDDREF pch l=0.04u w=0.12u
m19258 2995 3144 VDDREF VDDREF pch l=0.04u w=0.8u
m19259 VDDREF 3063 2996 VDDREF pch l=0.04u w=0.8u
m19260 2997 3146 VDDREF VDDREF pch l=0.04u w=0.8u
m19261 VDDREF 3064 2998 VDDREF pch l=0.04u w=0.8u
m19262 VDDREF 3206 2999 VDDREF pch l=0.04u w=0.8u
m19263 VDDREF 3207 3000 VDDREF pch l=0.04u w=0.8u
m19264 3001 3148 VDDREF VDDREF pch l=0.04u w=0.8u
m19265 VDDREF 3065 3002 VDDREF pch l=0.04u w=0.8u
m19266 VDDREF 131 3003 VDDREF pch l=0.04u w=0.8u
m19267 VDDREF 3066 3004 VDDREF pch l=0.04u w=0.8u
m19268 3005 3152 VDDREF VDDREF pch l=0.04u w=0.8u
m19269 VDDREF 3023 3006 VDDREF pch l=0.04u w=0.8u
m19270 VDDREF 3067 3007 VDDREF pch l=0.04u w=0.8u
m19271 VDDREF 3068 3008 VDDREF pch l=0.04u w=0.8u
m19272 3009 3156 VDDREF VDDREF pch l=0.04u w=0.8u
m19273 VDDREF 3024 3010 VDDREF pch l=0.04u w=0.8u
m19274 VDDREF FBDIV[9] 3011 VDDREF pch l=0.04u w=0.8u
m19275 VDDREF 3062 3012 VDDREF pch l=0.04u w=0.8u
m19276 3017 2955 VDDREF VDDREF pch l=0.04u w=0.8u
m19277 VDDREF 3041 3013 VDDREF pch l=0.04u w=0.8u
m19278 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19279 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19280 VDDREF 3015 3014 VDDREF pch l=0.04u w=1u
m19281 1146 2971 VDDREF VDDREF pch l=0.04u w=0.8u
m19282 3018 2972 VDDREF VDDREF pch l=0.04u w=0.8u
m19283 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19284 VDDREF 3023 30747 VDDREF pch l=0.04u w=0.12u
m19285 VDDREF 2796 30748 VDDREF pch l=0.04u w=0.12u
m19286 VDDREF 3024 30749 VDDREF pch l=0.04u w=0.12u
m19287 VDDREF 2799 30750 VDDREF pch l=0.04u w=0.12u
m19288 VDDREF 3044 2993 VDDREF pch l=0.04u w=0.8u
m19289 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19290 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19291 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19292 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19293 3019 2978 VDDREF VDDREF pch l=0.04u w=0.8u
m19294 3016 2508 2465 VDDREF pch l=0.04u w=0.8u
m19295 3020 437 VDDREF VDDREF pch l=0.04u w=0.8u
m19296 VDDREF 3046 2995 VDDREF pch l=0.04u w=0.8u
m19297 VDDREF 3048 2997 VDDREF pch l=0.04u w=0.8u
m19298 VDDREF 3050 3001 VDDREF pch l=0.04u w=0.8u
m19299 VDDREF 3055 3005 VDDREF pch l=0.04u w=0.8u
m19300 VDDREF 3059 3009 VDDREF pch l=0.04u w=0.8u
m19301 3012 3062 VDDREF VDDREF pch l=0.04u w=0.8u
m19302 3021 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19303 30760 3013 VDDREF VDDREF pch l=0.04u w=0.12u
m19304 3022 2970 VDDREF VDDREF pch l=0.04u w=0.8u
m19305 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19306 3023 2989 VDDREF VDDREF pch l=0.04u w=0.8u
m19307 2796 2990 VDDREF VDDREF pch l=0.04u w=0.8u
m19308 3024 2991 VDDREF VDDREF pch l=0.04u w=0.8u
m19309 2799 2992 VDDREF VDDREF pch l=0.04u w=0.8u
m19310 30762 2993 VDDREF VDDREF pch l=0.04u w=0.12u
m19311 2508 2465 3016 VDDREF pch l=0.04u w=0.8u
m19312 VDDREF 3062 3012 VDDREF pch l=0.04u w=0.8u
m19313 3026 3063 VDDREF VDDREF pch l=0.04u w=0.8u
m19314 3027 3064 VDDREF VDDREF pch l=0.04u w=0.8u
m19315 3028 2999 VDDREF VDDREF pch l=0.04u w=0.8u
m19316 3029 3000 VDDREF VDDREF pch l=0.04u w=0.8u
m19317 3030 3065 VDDREF VDDREF pch l=0.04u w=0.8u
m19318 3031 131 VDDREF VDDREF pch l=0.04u w=0.8u
m19319 3032 3066 VDDREF VDDREF pch l=0.04u w=0.8u
m19320 3033 3023 VDDREF VDDREF pch l=0.04u w=0.8u
m19321 3034 3067 VDDREF VDDREF pch l=0.04u w=0.8u
m19322 3035 3068 VDDREF VDDREF pch l=0.04u w=0.8u
m19323 3036 3024 VDDREF VDDREF pch l=0.04u w=0.8u
m19324 3037 FBDIV[9] VDDREF VDDREF pch l=0.04u w=0.8u
m19325 3039 3017 VDDREF VDDREF pch l=0.04u w=0.8u
m19326 3041 4251 30760 VDDREF pch l=0.04u w=0.12u
m19327 3040 3070 3022 VDDREF pch l=0.04u w=0.8u
m19328 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19329 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19330 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19331 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19332 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19333 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19334 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19335 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19336 3044 3085 30762 VDDREF pch l=0.04u w=0.12u
m19337 3042 912 VDDREF VDDREF pch l=0.04u w=0.8u
m19338 3043 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19339 3025 110 437 VDDREF pch l=0.04u w=0.8u
m19340 3046 2909 VDDREF VDDREF pch l=0.04u w=0.8u
m19341 3048 2911 VDDREF VDDREF pch l=0.04u w=0.8u
m19342 3050 2913 VDDREF VDDREF pch l=0.04u w=0.8u
m19343 3055 2917 VDDREF VDDREF pch l=0.04u w=0.8u
m19344 3059 2921 VDDREF VDDREF pch l=0.04u w=0.8u
m19345 3052 4328 3038 VDDREF pch l=0.04u w=0.8u
m19346 VDDREF 4351 3039 VDDREF pch l=0.04u w=0.8u
m19347 3069 3141 3041 VDDREF pch l=0.04u w=0.8u
m19348 3070 3022 3040 VDDREF pch l=0.04u w=0.8u
m19349 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19350 3071 4251 3044 VDDREF pch l=0.04u w=0.8u
m19351 3073 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19352 3074 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19353 3075 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19354 3076 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19355 3045 3016 VDDREF VDDREF pch l=0.04u w=0.8u
m19356 110 437 3025 VDDREF pch l=0.04u w=0.8u
m19357 VDDREF 2947 3046 VDDREF pch l=0.04u w=0.8u
m19358 VDDREF 2948 3048 VDDREF pch l=0.04u w=0.8u
m19359 VDDREF 2949 3050 VDDREF pch l=0.04u w=0.8u
m19360 VDDREF 2950 3055 VDDREF pch l=0.04u w=0.8u
m19361 VDDREF 2951 3059 VDDREF pch l=0.04u w=0.8u
m19362 VDDREF 4062 3062 VDDREF pch l=0.04u w=0.8u
m19363 3080 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19364 3081 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19365 3047 3065 3063 VDDREF pch l=0.04u w=0.8u
m19366 3049 1877 3064 VDDREF pch l=0.04u w=0.8u
m19367 3082 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19368 3083 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19369 3051 FRAC[9] 3065 VDDREF pch l=0.04u w=0.8u
m19370 30779 3021 3052 VDDREF pch l=0.04u w=0.12u
m19371 3053 3066 131 VDDREF pch l=0.04u w=0.8u
m19372 3054 3078 3066 VDDREF pch l=0.04u w=0.8u
m19373 3056 2900 3023 VDDREF pch l=0.04u w=0.8u
m19374 3057 2988 3067 VDDREF pch l=0.04u w=0.8u
m19375 3058 3079 3068 VDDREF pch l=0.04u w=0.8u
m19376 3060 FRAC[9] 3024 VDDREF pch l=0.04u w=0.8u
m19377 3061 2988 FBDIV[9] VDDREF pch l=0.04u w=0.8u
m19378 3039 3484 VDDREF VDDREF pch l=0.04u w=0.8u
m19379 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19380 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19381 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19382 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19383 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19384 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19385 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19386 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19387 3072 1146 912 VDDREF pch l=0.04u w=0.8u
m19388 3084 4328 3018 VDDREF pch l=0.04u w=0.8u
m19389 VDDREF 2844 3045 VDDREF pch l=0.04u w=0.8u
m19390 3065 3063 3047 VDDREF pch l=0.04u w=0.8u
m19391 1877 3064 3049 VDDREF pch l=0.04u w=0.8u
m19392 FRAC[9] 3065 3051 VDDREF pch l=0.04u w=0.8u
m19393 VDDREF 3101 30779 VDDREF pch l=0.04u w=0.12u
m19394 3066 131 3053 VDDREF pch l=0.04u w=0.8u
m19395 3078 3066 3054 VDDREF pch l=0.04u w=0.8u
m19396 2900 3023 3056 VDDREF pch l=0.04u w=0.8u
m19397 2988 3067 3057 VDDREF pch l=0.04u w=0.8u
m19398 3079 3068 3058 VDDREF pch l=0.04u w=0.8u
m19399 FRAC[9] 3024 3060 VDDREF pch l=0.04u w=0.8u
m19400 2988 FBDIV[9] 3061 VDDREF pch l=0.04u w=0.8u
m19401 VDDREF 3118 3069 VDDREF pch l=0.04u w=0.8u
m19402 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19403 VDDREF 4251 3085 VDDREF pch l=0.04u w=0.8u
m19404 1146 912 3072 VDDREF pch l=0.04u w=0.8u
m19405 30787 3043 3084 VDDREF pch l=0.04u w=0.12u
m19406 3092 4328 3086 VDDREF pch l=0.04u w=0.8u
m19407 3093 4328 2931 VDDREF pch l=0.04u w=0.8u
m19408 3094 4328 3087 VDDREF pch l=0.04u w=0.8u
m19409 3095 4328 2805 VDDREF pch l=0.04u w=0.8u
m19410 3096 3096 VDDREF VDDREF pch l=0.04u w=1u
m19411 3088 3025 VDDREF VDDREF pch l=0.04u w=0.8u
m19412 2947 2924 2925 VDDREF pch l=0.04u w=0.8u
m19413 2948 2930 2054 VDDREF pch l=0.04u w=0.8u
m19414 2949 2925 FRAC[15] VDDREF pch l=0.04u w=0.8u
m19415 3101 3052 VDDREF VDDREF pch l=0.04u w=0.8u
m19416 2950 2855 2745 VDDREF pch l=0.04u w=0.8u
m19417 2951 2857 FRAC[15] VDDREF pch l=0.04u w=0.8u
m19418 3102 3117 VDDREF VDDREF pch l=0.04u w=0.8u
m19419 3097 4328 3090 VDDREF pch l=0.04u w=0.8u
m19420 3098 4328 3091 VDDREF pch l=0.04u w=0.8u
m19421 3099 4328 3028 VDDREF pch l=0.04u w=0.8u
m19422 3100 4328 3029 VDDREF pch l=0.04u w=0.8u
m19423 3113 3039 VDDREF VDDREF pch l=0.04u w=0.8u
m19424 30792 3069 VDDREF VDDREF pch l=0.04u w=0.12u
m19425 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19426 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19427 3114 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m19428 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19429 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19430 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19431 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19432 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19433 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19434 VDDREF 3119 30787 VDDREF pch l=0.04u w=0.12u
m19435 30796 3073 3092 VDDREF pch l=0.04u w=0.12u
m19436 30797 3074 3093 VDDREF pch l=0.04u w=0.12u
m19437 30798 3075 3094 VDDREF pch l=0.04u w=0.12u
m19438 30799 3076 3095 VDDREF pch l=0.04u w=0.12u
m19439 3115 3045 VDDREF VDDREF pch l=0.04u w=0.8u
m19440 VDDREF 2860 3088 VDDREF pch l=0.04u w=0.8u
m19441 2924 2925 2947 VDDREF pch l=0.04u w=0.8u
m19442 2930 2054 2948 VDDREF pch l=0.04u w=0.8u
m19443 2925 FRAC[15] 2949 VDDREF pch l=0.04u w=0.8u
m19444 2855 2745 2950 VDDREF pch l=0.04u w=0.8u
m19445 2857 FRAC[15] 2951 VDDREF pch l=0.04u w=0.8u
m19446 3116 3122 3102 VDDREF pch l=0.04u w=0.8u
m19447 30804 3080 3097 VDDREF pch l=0.04u w=0.12u
m19448 30805 3081 3098 VDDREF pch l=0.04u w=0.12u
m19449 3103 3047 VDDREF VDDREF pch l=0.04u w=0.8u
m19450 3104 3049 VDDREF VDDREF pch l=0.04u w=0.8u
m19451 30806 3082 3099 VDDREF pch l=0.04u w=0.12u
m19452 30807 3083 3100 VDDREF pch l=0.04u w=0.12u
m19453 3105 3051 VDDREF VDDREF pch l=0.04u w=0.8u
m19454 3106 3053 VDDREF VDDREF pch l=0.04u w=0.8u
m19455 3107 3054 VDDREF VDDREF pch l=0.04u w=0.8u
m19456 3108 3056 VDDREF VDDREF pch l=0.04u w=0.8u
m19457 3109 3057 VDDREF VDDREF pch l=0.04u w=0.8u
m19458 3110 3058 VDDREF VDDREF pch l=0.04u w=0.8u
m19459 3111 3060 VDDREF VDDREF pch l=0.04u w=0.8u
m19460 3112 3061 VDDREF VDDREF pch l=0.04u w=0.8u
m19461 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19462 3118 3141 30792 VDDREF pch l=0.04u w=0.12u
m19463 3119 3084 VDDREF VDDREF pch l=0.04u w=0.8u
m19464 VDDREF 3132 30796 VDDREF pch l=0.04u w=0.12u
m19465 VDDREF 3133 30797 VDDREF pch l=0.04u w=0.12u
m19466 VDDREF 3134 30798 VDDREF pch l=0.04u w=0.12u
m19467 VDDREF 3135 30799 VDDREF pch l=0.04u w=0.12u
m19468 3071 3173 VDDREF VDDREF pch l=0.04u w=0.8u
m19469 2508 3120 VDDREF VDDREF pch l=0.04u w=0.8u
m19470 VDDREF 2946 3115 VDDREF pch l=0.04u w=0.8u
m19471 3122 3102 3116 VDDREF pch l=0.04u w=0.8u
m19472 VDDREF 3137 30804 VDDREF pch l=0.04u w=0.12u
m19473 VDDREF 3138 30805 VDDREF pch l=0.04u w=0.12u
m19474 VDDREF 2869 3103 VDDREF pch l=0.04u w=0.8u
m19475 VDDREF 2870 3104 VDDREF pch l=0.04u w=0.8u
m19476 VDDREF 3139 30806 VDDREF pch l=0.04u w=0.12u
m19477 VDDREF 3140 30807 VDDREF pch l=0.04u w=0.12u
m19478 VDDREF 2871 3105 VDDREF pch l=0.04u w=0.8u
m19479 3121 3021 3101 VDDREF pch l=0.04u w=0.8u
m19480 VDDREF 2872 3106 VDDREF pch l=0.04u w=0.8u
m19481 VDDREF 2873 3107 VDDREF pch l=0.04u w=0.8u
m19482 VDDREF 2874 3108 VDDREF pch l=0.04u w=0.8u
m19483 VDDREF 2875 3109 VDDREF pch l=0.04u w=0.8u
m19484 VDDREF 2876 3110 VDDREF pch l=0.04u w=0.8u
m19485 VDDREF 2877 3111 VDDREF pch l=0.04u w=0.8u
m19486 VDDREF 2878 3112 VDDREF pch l=0.04u w=0.8u
m19487 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19488 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19489 3128 4251 3118 VDDREF pch l=0.04u w=0.8u
m19490 3129 3113 VDDREF VDDREF pch l=0.04u w=0.8u
m19491 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19492 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19493 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19494 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19495 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19496 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19497 3130 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m19498 3131 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19499 3132 3092 VDDREF VDDREF pch l=0.04u w=0.8u
m19500 3133 3093 VDDREF VDDREF pch l=0.04u w=0.8u
m19501 3134 3094 VDDREF VDDREF pch l=0.04u w=0.8u
m19502 3135 3095 VDDREF VDDREF pch l=0.04u w=0.8u
m19503 VDDREF 3218 3071 VDDREF pch l=0.04u w=0.8u
m19504 3136 3088 VDDREF VDDREF pch l=0.04u w=0.8u
m19505 3137 3097 VDDREF VDDREF pch l=0.04u w=0.8u
m19506 3138 3098 VDDREF VDDREF pch l=0.04u w=0.8u
m19507 VDDREF 2924 3123 VDDREF pch l=0.04u w=0.8u
m19508 VDDREF 2930 3124 VDDREF pch l=0.04u w=0.8u
m19509 3139 3099 VDDREF VDDREF pch l=0.04u w=0.8u
m19510 3140 3100 VDDREF VDDREF pch l=0.04u w=0.8u
m19511 VDDREF 2925 3125 VDDREF pch l=0.04u w=0.8u
m19512 30816 4328 3121 VDDREF pch l=0.04u w=0.12u
m19513 VDDREF 2855 3126 VDDREF pch l=0.04u w=0.8u
m19514 VDDREF 2857 3127 VDDREF pch l=0.04u w=0.8u
m19515 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19516 VDDREF 3953 3129 VDDREF pch l=0.04u w=0.8u
m19517 VDDREF 1962 3130 VDDREF pch l=0.04u w=0.8u
m19518 3071 3218 VDDREF VDDREF pch l=0.04u w=0.8u
m19519 3142 3043 3119 VDDREF pch l=0.04u w=0.8u
m19520 3143 3016 VDDREF VDDREF pch l=0.04u w=0.8u
m19521 VDDREF 2979 3136 VDDREF pch l=0.04u w=0.8u
m19522 VDDREF 3169 30816 VDDREF pch l=0.04u w=0.12u
m19523 3145 3103 VDDREF VDDREF pch l=0.04u w=0.8u
m19524 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19525 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19526 3147 3104 VDDREF VDDREF pch l=0.04u w=0.8u
m19527 3149 3105 VDDREF VDDREF pch l=0.04u w=0.8u
m19528 3150 3106 VDDREF VDDREF pch l=0.04u w=0.8u
m19529 3151 3107 VDDREF VDDREF pch l=0.04u w=0.8u
m19530 3153 3108 VDDREF VDDREF pch l=0.04u w=0.8u
m19531 3154 3109 VDDREF VDDREF pch l=0.04u w=0.8u
m19532 3155 3110 VDDREF VDDREF pch l=0.04u w=0.8u
m19533 3157 3111 VDDREF VDDREF pch l=0.04u w=0.8u
m19534 3158 3112 VDDREF VDDREF pch l=0.04u w=0.8u
m19535 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19536 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19537 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19538 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19539 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19540 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19541 VDDREF 4251 3141 VDDREF pch l=0.04u w=0.8u
m19542 3159 4328 3072 VDDREF pch l=0.04u w=0.8u
m19543 VDDREF 3173 3071 VDDREF pch l=0.04u w=0.8u
m19544 30830 4328 3142 VDDREF pch l=0.04u w=0.12u
m19545 3160 3073 3132 VDDREF pch l=0.04u w=0.8u
m19546 3161 3074 3133 VDDREF pch l=0.04u w=0.8u
m19547 3162 3075 3134 VDDREF pch l=0.04u w=0.8u
m19548 3163 3076 3135 VDDREF pch l=0.04u w=0.8u
m19549 VDDREF 3174 VDDREF VDDREF pch l=0.26u w=1u
m19550 3169 3121 VDDREF VDDREF pch l=0.04u w=0.8u
m19551 3165 3080 3137 VDDREF pch l=0.04u w=0.8u
m19552 3166 3081 3138 VDDREF pch l=0.04u w=0.8u
m19553 3144 2924 VDDREF VDDREF pch l=0.04u w=0.8u
m19554 VDDREF 2996 3145 VDDREF pch l=0.04u w=0.8u
m19555 3146 2930 VDDREF VDDREF pch l=0.04u w=0.8u
m19556 VDDREF 2998 3147 VDDREF pch l=0.04u w=0.8u
m19557 3167 3082 3139 VDDREF pch l=0.04u w=0.8u
m19558 3168 3083 3140 VDDREF pch l=0.04u w=0.8u
m19559 3148 2925 VDDREF VDDREF pch l=0.04u w=0.8u
m19560 VDDREF 3002 3149 VDDREF pch l=0.04u w=0.8u
m19561 VDDREF 3003 3150 VDDREF pch l=0.04u w=0.8u
m19562 VDDREF 3004 3151 VDDREF pch l=0.04u w=0.8u
m19563 3152 2855 VDDREF VDDREF pch l=0.04u w=0.8u
m19564 VDDREF 3006 3153 VDDREF pch l=0.04u w=0.8u
m19565 VDDREF 3007 3154 VDDREF pch l=0.04u w=0.8u
m19566 VDDREF 3008 3155 VDDREF pch l=0.04u w=0.8u
m19567 3156 2857 VDDREF VDDREF pch l=0.04u w=0.8u
m19568 VDDREF 3010 3157 VDDREF pch l=0.04u w=0.8u
m19569 VDDREF 3011 3158 VDDREF pch l=0.04u w=0.8u
m19570 3170 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m19571 3171 3129 VDDREF VDDREF pch l=0.04u w=0.8u
m19572 3172 3114 VDDREF VDDREF pch l=0.04u w=0.8u
m19573 30834 3131 3159 VDDREF pch l=0.04u w=0.12u
m19574 VDDREF 61 30830 VDDREF pch l=0.04u w=0.12u
m19575 30837 4328 3160 VDDREF pch l=0.04u w=0.12u
m19576 30838 4328 3161 VDDREF pch l=0.04u w=0.12u
m19577 30839 4328 3162 VDDREF pch l=0.04u w=0.12u
m19578 30840 4328 3163 VDDREF pch l=0.04u w=0.12u
m19579 3175 3175 VDDREF VDDREF pch l=0.04u w=1u
m19580 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19581 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19582 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19583 3164 2844 3016 VDDREF pch l=0.04u w=0.8u
m19584 3176 3025 VDDREF VDDREF pch l=0.04u w=0.8u
m19585 30841 4328 3165 VDDREF pch l=0.04u w=0.12u
m19586 30842 4328 3166 VDDREF pch l=0.04u w=0.12u
m19587 VDDREF 2925 3144 VDDREF pch l=0.04u w=0.8u
m19588 VDDREF 2054 3146 VDDREF pch l=0.04u w=0.8u
m19589 30843 4328 3167 VDDREF pch l=0.04u w=0.12u
m19590 30844 4328 3168 VDDREF pch l=0.04u w=0.12u
m19591 VDDREF FRAC[15] 3148 VDDREF pch l=0.04u w=0.8u
m19592 VDDREF 3182 VDDREF VDDREF pch l=0.26u w=1u
m19593 VDDREF 2745 3152 VDDREF pch l=0.04u w=0.8u
m19594 VDDREF FRAC[15] 3156 VDDREF pch l=0.04u w=0.8u
m19595 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19596 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19597 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19598 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19599 3177 3199 3171 VDDREF pch l=0.04u w=0.8u
m19600 3128 3249 VDDREF VDDREF pch l=0.04u w=0.8u
m19601 VDDREF 3040 3172 VDDREF pch l=0.04u w=0.8u
m19602 VDDREF 3200 30834 VDDREF pch l=0.04u w=0.12u
m19603 61 3142 VDDREF VDDREF pch l=0.04u w=0.8u
m19604 VDDREF 3201 30837 VDDREF pch l=0.04u w=0.12u
m19605 VDDREF 2797 30838 VDDREF pch l=0.04u w=0.12u
m19606 VDDREF 3202 30839 VDDREF pch l=0.04u w=0.12u
m19607 VDDREF 2800 30840 VDDREF pch l=0.04u w=0.12u
m19608 3173 3301 VDDREF VDDREF pch l=0.04u w=0.8u
m19609 2844 3016 3164 VDDREF pch l=0.04u w=0.8u
m19610 VDDREF 3203 30841 VDDREF pch l=0.04u w=0.12u
m19611 VDDREF 3063 30842 VDDREF pch l=0.04u w=0.12u
m19612 VDDREF 3204 30843 VDDREF pch l=0.04u w=0.12u
m19613 VDDREF 3065 30844 VDDREF pch l=0.04u w=0.12u
m19614 3181 3181 VDDREF VDDREF pch l=0.04u w=1u
m19615 3184 3047 VDDREF VDDREF pch l=0.04u w=0.8u
m19616 3186 3049 VDDREF VDDREF pch l=0.04u w=0.8u
m19617 3188 3051 VDDREF VDDREF pch l=0.04u w=0.8u
m19618 3189 3053 VDDREF VDDREF pch l=0.04u w=0.8u
m19619 3190 3054 VDDREF VDDREF pch l=0.04u w=0.8u
m19620 3192 3056 VDDREF VDDREF pch l=0.04u w=0.8u
m19621 3193 3057 VDDREF VDDREF pch l=0.04u w=0.8u
m19622 3194 3058 VDDREF VDDREF pch l=0.04u w=0.8u
m19623 3196 3060 VDDREF VDDREF pch l=0.04u w=0.8u
m19624 3197 3061 VDDREF VDDREF pch l=0.04u w=0.8u
m19625 3198 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m19626 3199 3171 3177 VDDREF pch l=0.04u w=0.8u
m19627 VDDREF 3290 3128 VDDREF pch l=0.04u w=0.8u
m19628 3200 3159 VDDREF VDDREF pch l=0.04u w=0.8u
m19629 3201 3160 VDDREF VDDREF pch l=0.04u w=0.8u
m19630 2797 3161 VDDREF VDDREF pch l=0.04u w=0.8u
m19631 3202 3162 VDDREF VDDREF pch l=0.04u w=0.8u
m19632 2800 3163 VDDREF VDDREF pch l=0.04u w=0.8u
m19633 VDDREF 3272 3173 VDDREF pch l=0.04u w=0.8u
m19634 VDDREF 3213 VDDREF VDDREF pch l=0.26u w=1u
m19635 VDDREF 3216 VDDREF VDDREF pch l=0.26u w=1u
m19636 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19637 VDDREF 3178 3179 VDDREF pch l=0.04u w=1u
m19638 3203 3165 VDDREF VDDREF pch l=0.04u w=0.8u
m19639 3063 3166 VDDREF VDDREF pch l=0.04u w=0.8u
m19640 VDDREF 3219 VDDREF VDDREF pch l=0.26u w=1u
m19641 VDDREF 3222 VDDREF VDDREF pch l=0.26u w=1u
m19642 3204 3167 VDDREF VDDREF pch l=0.04u w=0.8u
m19643 3065 3168 VDDREF VDDREF pch l=0.04u w=0.8u
m19644 VDDREF 3223 VDDREF VDDREF pch l=0.26u w=1u
m19645 VDDREF 3226 VDDREF VDDREF pch l=0.26u w=1u
m19646 30855 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m19647 3180 2860 3025 VDDREF pch l=0.04u w=0.8u
m19648 3090 3228 3183 VDDREF pch l=0.04u w=0.8u
m19649 3206 3229 3185 VDDREF pch l=0.04u w=0.8u
m19650 3208 3230 3187 VDDREF pch l=0.04u w=0.8u
m19651 2742 3231 3191 VDDREF pch l=0.04u w=0.8u
m19652 2744 3232 3195 VDDREF pch l=0.04u w=0.8u
m19653 VDDREF 320 3198 VDDREF pch l=0.04u w=0.8u
m19654 3128 3290 VDDREF VDDREF pch l=0.04u w=0.8u
m19655 3212 3172 VDDREF VDDREF pch l=0.04u w=0.8u
m19656 3214 3214 VDDREF VDDREF pch l=0.04u w=1u
m19657 3215 3215 VDDREF VDDREF pch l=0.04u w=1u
m19658 3217 2098 VDDREF VDDREF pch l=0.04u w=0.8u
m19659 3220 3220 VDDREF VDDREF pch l=0.04u w=1u
m19660 3221 3221 VDDREF VDDREF pch l=0.04u w=1u
m19661 3224 3224 VDDREF VDDREF pch l=0.04u w=1u
m19662 3225 3225 VDDREF VDDREF pch l=0.04u w=1u
m19663 3205 3164 30855 VDDREF pch l=0.04u w=0.8u
m19664 3227 2508 VDDREF VDDREF pch l=0.04u w=0.8u
m19665 2860 3025 3180 VDDREF pch l=0.04u w=0.8u
m19666 3228 3183 3090 VDDREF pch l=0.04u w=0.8u
m19667 3229 3185 3206 VDDREF pch l=0.04u w=0.8u
m19668 3230 3187 3208 VDDREF pch l=0.04u w=0.8u
m19669 VDDREF 3210 3209 VDDREF pch l=0.04u w=1u
m19670 3231 3191 2742 VDDREF pch l=0.04u w=0.8u
m19671 3232 3195 2744 VDDREF pch l=0.04u w=0.8u
m19672 3091 2869 3047 VDDREF pch l=0.04u w=0.8u
m19673 3207 2870 3049 VDDREF pch l=0.04u w=0.8u
m19674 3064 2871 3051 VDDREF pch l=0.04u w=0.8u
m19675 3038 2872 3053 VDDREF pch l=0.04u w=0.8u
m19676 3211 2873 3054 VDDREF pch l=0.04u w=0.8u
m19677 2898 2874 3056 VDDREF pch l=0.04u w=0.8u
m19678 3078 2875 3057 VDDREF pch l=0.04u w=0.8u
m19679 3067 2876 3058 VDDREF pch l=0.04u w=0.8u
m19680 2900 2877 3060 VDDREF pch l=0.04u w=0.8u
m19681 3079 2878 3061 VDDREF pch l=0.04u w=0.8u
m19682 VDDREF 3249 3128 VDDREF pch l=0.04u w=0.8u
m19683 VDDREF 3130 3212 VDDREF pch l=0.04u w=0.8u
m19684 3233 3131 3200 VDDREF pch l=0.04u w=0.8u
m19685 VDDREF 3252 VDDREF VDDREF pch l=0.26u w=1u
m19686 3235 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19687 3236 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19688 3237 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19689 3238 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19690 3218 FBDIV[10] VDDREF VDDREF pch l=0.04u w=0.8u
m19691 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m19692 VDDREF 2906 3227 VDDREF pch l=0.04u w=0.8u
m19693 2869 3047 3091 VDDREF pch l=0.04u w=0.8u
m19694 2870 3049 3207 VDDREF pch l=0.04u w=0.8u
m19695 2871 3051 3064 VDDREF pch l=0.04u w=0.8u
m19696 2872 3053 3038 VDDREF pch l=0.04u w=0.8u
m19697 2873 3054 3211 VDDREF pch l=0.04u w=0.8u
m19698 2874 3056 2898 VDDREF pch l=0.04u w=0.8u
m19699 2875 3057 3078 VDDREF pch l=0.04u w=0.8u
m19700 2876 3058 3067 VDDREF pch l=0.04u w=0.8u
m19701 2877 3060 2900 VDDREF pch l=0.04u w=0.8u
m19702 2878 3061 3079 VDDREF pch l=0.04u w=0.8u
m19703 3248 3170 VDDREF VDDREF pch l=0.04u w=0.8u
m19704 3250 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m19705 3212 3130 VDDREF VDDREF pch l=0.04u w=0.8u
m19706 30884 4328 3233 VDDREF pch l=0.04u w=0.12u
m19707 3251 3251 VDDREF VDDREF pch l=0.04u w=1u
m19708 VDDREF 4062 3218 VDDREF pch l=0.04u w=0.8u
m19709 VDDREF 3239 3240 VDDREF pch l=0.04u w=1u
m19710 VDDREF 3242 3241 VDDREF pch l=0.04u w=1u
m19711 3234 3018 2098 VDDREF pch l=0.04u w=0.8u
m19712 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m19713 3255 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m19714 3256 110 VDDREF VDDREF pch l=0.04u w=0.8u
m19715 VDDREF 3228 3243 VDDREF pch l=0.04u w=0.8u
m19716 VDDREF 3229 3244 VDDREF pch l=0.04u w=0.8u
m19717 VDDREF 3230 3245 VDDREF pch l=0.04u w=0.8u
m19718 VDDREF 3231 3246 VDDREF pch l=0.04u w=0.8u
m19719 VDDREF 3232 3247 VDDREF pch l=0.04u w=0.8u
m19720 VDDREF 3116 3248 VDDREF pch l=0.04u w=0.8u
m19721 3249 3381 VDDREF VDDREF pch l=0.04u w=0.8u
m19722 VDDREF 3172 3212 VDDREF pch l=0.04u w=0.8u
m19723 VDDREF 3287 30884 VDDREF pch l=0.04u w=0.12u
m19724 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m19725 3018 2098 3234 VDDREF pch l=0.04u w=0.8u
m19726 3266 4328 3253 VDDREF pch l=0.04u w=0.8u
m19727 3267 4328 3211 VDDREF pch l=0.04u w=0.8u
m19728 3268 4328 3254 VDDREF pch l=0.04u w=0.8u
m19729 3269 4328 3067 VDDREF pch l=0.04u w=0.8u
m19730 VDDREF 2906 3255 VDDREF pch l=0.04u w=0.8u
m19731 3273 2906 VDDREF VDDREF pch l=0.04u w=0.8u
m19732 VDDREF 731 3256 VDDREF pch l=0.04u w=0.8u
m19733 VDDREF 3257 3258 VDDREF pch l=0.04u w=1u
m19734 VDDREF 3260 3259 VDDREF pch l=0.04u w=1u
m19735 3274 3338 VDDREF VDDREF pch l=0.04u w=0.8u
m19736 3275 1908 VDDREF VDDREF pch l=0.04u w=0.8u
m19737 3276 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m19738 3277 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m19739 VDDREF 3261 3262 VDDREF pch l=0.04u w=1u
m19740 VDDREF 3264 3263 VDDREF pch l=0.04u w=1u
m19741 3278 FRAC[10] VDDREF VDDREF pch l=0.04u w=0.8u
m19742 VDDREF 3315 3265 VDDREF pch l=0.04u w=0.8u
m19743 3279 3339 VDDREF VDDREF pch l=0.04u w=0.8u
m19744 3280 3352 VDDREF VDDREF pch l=0.04u w=0.8u
m19745 3281 3254 VDDREF VDDREF pch l=0.04u w=0.8u
m19746 3282 3265 VDDREF VDDREF pch l=0.04u w=0.8u
m19747 3283 3353 VDDREF VDDREF pch l=0.04u w=0.8u
m19748 3284 FRAC[10] VDDREF VDDREF pch l=0.04u w=0.8u
m19749 3285 3265 VDDREF VDDREF pch l=0.04u w=0.8u
m19750 VDDREF 3344 3249 VDDREF pch l=0.04u w=0.8u
m19751 3286 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m19752 3287 3233 VDDREF VDDREF pch l=0.04u w=0.8u
m19753 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m19754 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m19755 VDDREF 3271 3270 VDDREF pch l=0.04u w=1u
m19756 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m19757 30903 3235 3266 VDDREF pch l=0.04u w=0.12u
m19758 30904 3236 3267 VDDREF pch l=0.04u w=0.12u
m19759 30905 3237 3268 VDDREF pch l=0.04u w=0.12u
m19760 30906 3238 3269 VDDREF pch l=0.04u w=0.12u
m19761 VDDREF 4062 3272 VDDREF pch l=0.04u w=0.8u
m19762 2909 3412 VDDREF VDDREF pch l=0.04u w=0.8u
m19763 VDDREF 3336 3274 VDDREF pch l=0.04u w=0.8u
m19764 2911 3414 VDDREF VDDREF pch l=0.04u w=0.8u
m19765 VDDREF 3337 3275 VDDREF pch l=0.04u w=0.8u
m19766 VDDREF 3481 3276 VDDREF pch l=0.04u w=0.8u
m19767 VDDREF 3482 3277 VDDREF pch l=0.04u w=0.8u
m19768 2913 3416 VDDREF VDDREF pch l=0.04u w=0.8u
m19769 VDDREF 3338 3278 VDDREF pch l=0.04u w=0.8u
m19770 VDDREF 131 3279 VDDREF pch l=0.04u w=0.8u
m19771 VDDREF 3339 3280 VDDREF pch l=0.04u w=0.8u
m19772 2917 3420 VDDREF VDDREF pch l=0.04u w=0.8u
m19773 VDDREF 3340 3281 VDDREF pch l=0.04u w=0.8u
m19774 VDDREF 3341 3282 VDDREF pch l=0.04u w=0.8u
m19775 VDDREF 3342 3283 VDDREF pch l=0.04u w=0.8u
m19776 2921 3424 VDDREF VDDREF pch l=0.04u w=0.8u
m19777 VDDREF 3343 3284 VDDREF pch l=0.04u w=0.8u
m19778 VDDREF FBDIV[10] 3285 VDDREF pch l=0.04u w=0.8u
m19779 3289 3248 VDDREF VDDREF pch l=0.04u w=0.8u
m19780 VDDREF FBDIV[11] 3286 VDDREF pch l=0.04u w=0.8u
m19781 3291 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m19782 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m19783 VDDREF 3297 30903 VDDREF pch l=0.04u w=0.12u
m19784 VDDREF 3298 30904 VDDREF pch l=0.04u w=0.12u
m19785 VDDREF 3299 30905 VDDREF pch l=0.04u w=0.12u
m19786 VDDREF 3300 30906 VDDREF pch l=0.04u w=0.12u
m19787 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m19788 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m19789 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m19790 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m19791 3293 3255 VDDREF VDDREF pch l=0.04u w=0.8u
m19792 3288 2508 2906 VDDREF pch l=0.04u w=0.8u
m19793 3294 731 VDDREF VDDREF pch l=0.04u w=0.8u
m19794 VDDREF 3320 2909 VDDREF pch l=0.04u w=0.8u
m19795 VDDREF 3322 2911 VDDREF pch l=0.04u w=0.8u
m19796 VDDREF 3324 2913 VDDREF pch l=0.04u w=0.8u
m19797 VDDREF 3329 2917 VDDREF pch l=0.04u w=0.8u
m19798 VDDREF 3333 2921 VDDREF pch l=0.04u w=0.8u
m19799 VDDREF 3198 3289 VDDREF pch l=0.04u w=0.8u
m19800 3295 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19801 3290 1676 VDDREF VDDREF pch l=0.04u w=0.8u
m19802 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m19803 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m19804 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m19805 VDDREF 3287 3292 VDDREF pch l=0.04u w=0.8u
m19806 3296 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19807 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m19808 3297 3266 VDDREF VDDREF pch l=0.04u w=0.8u
m19809 3298 3267 VDDREF VDDREF pch l=0.04u w=0.8u
m19810 3299 3268 VDDREF VDDREF pch l=0.04u w=0.8u
m19811 3300 3269 VDDREF VDDREF pch l=0.04u w=0.8u
m19812 2508 2906 3288 VDDREF pch l=0.04u w=0.8u
m19813 3289 3198 VDDREF VDDREF pch l=0.04u w=0.8u
m19814 3303 3336 VDDREF VDDREF pch l=0.04u w=0.8u
m19815 3304 3337 VDDREF VDDREF pch l=0.04u w=0.8u
m19816 3305 3276 VDDREF VDDREF pch l=0.04u w=0.8u
m19817 3306 3277 VDDREF VDDREF pch l=0.04u w=0.8u
m19818 3307 3338 VDDREF VDDREF pch l=0.04u w=0.8u
m19819 3308 131 VDDREF VDDREF pch l=0.04u w=0.8u
m19820 3309 3339 VDDREF VDDREF pch l=0.04u w=0.8u
m19821 3310 3340 VDDREF VDDREF pch l=0.04u w=0.8u
m19822 3311 3341 VDDREF VDDREF pch l=0.04u w=0.8u
m19823 3312 3342 VDDREF VDDREF pch l=0.04u w=0.8u
m19824 3313 3343 VDDREF VDDREF pch l=0.04u w=0.8u
m19825 3314 FBDIV[10] VDDREF VDDREF pch l=0.04u w=0.8u
m19826 VDDREF 4062 3290 VDDREF pch l=0.04u w=0.8u
m19827 3317 3250 VDDREF VDDREF pch l=0.04u w=0.8u
m19828 3316 4251 3212 VDDREF pch l=0.04u w=0.8u
m19829 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m19830 415 3292 VDDREF VDDREF pch l=0.04u w=0.8u
m19831 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m19832 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m19833 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m19834 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m19835 3301 3350 2926 VDDREF pch l=0.04u w=0.8u
m19836 VDDREF 3248 3289 VDDREF pch l=0.04u w=0.8u
m19837 3302 110 731 VDDREF pch l=0.04u w=0.8u
m19838 3320 3183 VDDREF VDDREF pch l=0.04u w=0.8u
m19839 3322 3185 VDDREF VDDREF pch l=0.04u w=0.8u
m19840 3324 3187 VDDREF VDDREF pch l=0.04u w=0.8u
m19841 3329 3191 VDDREF VDDREF pch l=0.04u w=0.8u
m19842 3333 3195 VDDREF VDDREF pch l=0.04u w=0.8u
m19843 3326 4328 3315 VDDREF pch l=0.04u w=0.8u
m19844 VDDREF 3177 3317 VDDREF pch l=0.04u w=0.8u
m19845 30928 3291 3316 VDDREF pch l=0.04u w=0.12u
m19846 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m19847 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m19848 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m19849 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m19850 3345 4328 3234 VDDREF pch l=0.04u w=0.8u
m19851 3346 3235 3297 VDDREF pch l=0.04u w=0.8u
m19852 3347 3236 3298 VDDREF pch l=0.04u w=0.8u
m19853 3348 3237 3299 VDDREF pch l=0.04u w=0.8u
m19854 3349 3238 3300 VDDREF pch l=0.04u w=0.8u
m19855 3350 2926 3301 VDDREF pch l=0.04u w=0.8u
m19856 3319 3288 VDDREF VDDREF pch l=0.04u w=0.8u
m19857 110 731 3302 VDDREF pch l=0.04u w=0.8u
m19858 VDDREF 3228 3320 VDDREF pch l=0.04u w=0.8u
m19859 VDDREF 3229 3322 VDDREF pch l=0.04u w=0.8u
m19860 VDDREF 3230 3324 VDDREF pch l=0.04u w=0.8u
m19861 VDDREF 3231 3329 VDDREF pch l=0.04u w=0.8u
m19862 VDDREF 3232 3333 VDDREF pch l=0.04u w=0.8u
m19863 3354 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19864 3355 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19865 3321 3338 3336 VDDREF pch l=0.04u w=0.8u
m19866 3323 1908 3337 VDDREF pch l=0.04u w=0.8u
m19867 3356 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19868 3357 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19869 3325 FRAC[10] 3338 VDDREF pch l=0.04u w=0.8u
m19870 30933 3295 3326 VDDREF pch l=0.04u w=0.12u
m19871 3327 3339 131 VDDREF pch l=0.04u w=0.8u
m19872 3328 3352 3339 VDDREF pch l=0.04u w=0.8u
m19873 3330 3254 3340 VDDREF pch l=0.04u w=0.8u
m19874 3331 3265 3341 VDDREF pch l=0.04u w=0.8u
m19875 3332 3353 3342 VDDREF pch l=0.04u w=0.8u
m19876 3334 FRAC[10] 3343 VDDREF pch l=0.04u w=0.8u
m19877 3335 3265 FBDIV[10] VDDREF pch l=0.04u w=0.8u
m19878 VDDREF 4062 3344 VDDREF pch l=0.04u w=0.8u
m19879 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m19880 VDDREF 3364 30928 VDDREF pch l=0.04u w=0.12u
m19881 3358 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19882 30940 3296 3345 VDDREF pch l=0.04u w=0.12u
m19883 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m19884 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m19885 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m19886 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m19887 30941 4328 3346 VDDREF pch l=0.04u w=0.12u
m19888 30942 4328 3347 VDDREF pch l=0.04u w=0.12u
m19889 30943 4328 3348 VDDREF pch l=0.04u w=0.12u
m19890 30944 4328 3349 VDDREF pch l=0.04u w=0.12u
m19891 VDDREF 3318 3350 VDDREF pch l=0.04u w=0.8u
m19892 VDDREF 3115 3319 VDDREF pch l=0.04u w=0.8u
m19893 3359 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m19894 3338 3336 3321 VDDREF pch l=0.04u w=0.8u
m19895 1908 3337 3323 VDDREF pch l=0.04u w=0.8u
m19896 FRAC[10] 3338 3325 VDDREF pch l=0.04u w=0.8u
m19897 VDDREF 3370 30933 VDDREF pch l=0.04u w=0.12u
m19898 3339 131 3327 VDDREF pch l=0.04u w=0.8u
m19899 3352 3339 3328 VDDREF pch l=0.04u w=0.8u
m19900 3254 3340 3330 VDDREF pch l=0.04u w=0.8u
m19901 3265 3341 3331 VDDREF pch l=0.04u w=0.8u
m19902 3353 3342 3332 VDDREF pch l=0.04u w=0.8u
m19903 FRAC[10] 3343 3334 VDDREF pch l=0.04u w=0.8u
m19904 3265 FBDIV[10] 3335 VDDREF pch l=0.04u w=0.8u
m19905 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m19906 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m19907 3364 3316 VDDREF VDDREF pch l=0.04u w=0.8u
m19908 3365 3317 VDDREF VDDREF pch l=0.04u w=0.8u
m19909 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m19910 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m19911 VDDREF 3383 30940 VDDREF pch l=0.04u w=0.12u
m19912 VDDREF 3340 30941 VDDREF pch l=0.04u w=0.12u
m19913 VDDREF 3066 30942 VDDREF pch l=0.04u w=0.12u
m19914 VDDREF 3343 30943 VDDREF pch l=0.04u w=0.12u
m19915 VDDREF 3068 30944 VDDREF pch l=0.04u w=0.12u
m19916 3360 3302 VDDREF VDDREF pch l=0.04u w=0.8u
m19917 3228 3203 3204 VDDREF pch l=0.04u w=0.8u
m19918 3229 3208 2024 VDDREF pch l=0.04u w=0.8u
m19919 3230 3204 FRAC[14] VDDREF pch l=0.04u w=0.8u
m19920 3370 3326 VDDREF VDDREF pch l=0.04u w=0.8u
m19921 3231 2854 2744 VDDREF pch l=0.04u w=0.8u
m19922 3232 2856 FRAC[14] VDDREF pch l=0.04u w=0.8u
m19923 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m19924 3366 4328 3362 VDDREF pch l=0.04u w=0.8u
m19925 3367 4328 3363 VDDREF pch l=0.04u w=0.8u
m19926 3368 4328 3305 VDDREF pch l=0.04u w=0.8u
m19927 3369 4328 3306 VDDREF pch l=0.04u w=0.8u
m19928 VDDREF 3286 3365 VDDREF pch l=0.04u w=0.8u
m19929 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m19930 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m19931 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m19932 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m19933 3383 3345 VDDREF VDDREF pch l=0.04u w=0.8u
m19934 3382 4328 3287 VDDREF pch l=0.04u w=0.8u
m19935 3340 3346 VDDREF VDDREF pch l=0.04u w=0.8u
m19936 3066 3347 VDDREF VDDREF pch l=0.04u w=0.8u
m19937 3343 3348 VDDREF VDDREF pch l=0.04u w=0.8u
m19938 3068 3349 VDDREF VDDREF pch l=0.04u w=0.8u
m19939 3318 3953 VDDREF VDDREF pch l=0.04u w=0.8u
m19940 3385 3319 VDDREF VDDREF pch l=0.04u w=0.8u
m19941 VDDREF 3136 3360 VDDREF pch l=0.04u w=0.8u
m19942 3203 3204 3228 VDDREF pch l=0.04u w=0.8u
m19943 3208 2024 3229 VDDREF pch l=0.04u w=0.8u
m19944 3204 FRAC[14] 3230 VDDREF pch l=0.04u w=0.8u
m19945 2854 2744 3231 VDDREF pch l=0.04u w=0.8u
m19946 2856 FRAC[14] 3232 VDDREF pch l=0.04u w=0.8u
m19947 3384 4251 3289 VDDREF pch l=0.04u w=0.8u
m19948 30959 3354 3366 VDDREF pch l=0.04u w=0.12u
m19949 30960 3355 3367 VDDREF pch l=0.04u w=0.12u
m19950 3371 3321 VDDREF VDDREF pch l=0.04u w=0.8u
m19951 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m19952 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m19953 3372 3323 VDDREF VDDREF pch l=0.04u w=0.8u
m19954 30961 3356 3368 VDDREF pch l=0.04u w=0.12u
m19955 30962 3357 3369 VDDREF pch l=0.04u w=0.12u
m19956 3373 3325 VDDREF VDDREF pch l=0.04u w=0.8u
m19957 3374 3327 VDDREF VDDREF pch l=0.04u w=0.8u
m19958 3375 3328 VDDREF VDDREF pch l=0.04u w=0.8u
m19959 3376 3330 VDDREF VDDREF pch l=0.04u w=0.8u
m19960 3377 3331 VDDREF VDDREF pch l=0.04u w=0.8u
m19961 3378 3332 VDDREF VDDREF pch l=0.04u w=0.8u
m19962 3379 3334 VDDREF VDDREF pch l=0.04u w=0.8u
m19963 3380 3335 VDDREF VDDREF pch l=0.04u w=0.8u
m19964 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m19965 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m19966 3365 3286 VDDREF VDDREF pch l=0.04u w=0.8u
m19967 3381 3394 3013 VDDREF pch l=0.04u w=0.8u
m19968 3387 3291 3364 VDDREF pch l=0.04u w=0.8u
m19969 30969 3358 3382 VDDREF pch l=0.04u w=0.12u
m19970 VDDREF 3400 3318 VDDREF pch l=0.04u w=0.8u
m19971 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m19972 VDDREF 3227 3385 VDDREF pch l=0.04u w=0.8u
m19973 30972 3359 3384 VDDREF pch l=0.04u w=0.12u
m19974 VDDREF 3402 30959 VDDREF pch l=0.04u w=0.12u
m19975 VDDREF 3403 30960 VDDREF pch l=0.04u w=0.12u
m19976 VDDREF 3145 3371 VDDREF pch l=0.04u w=0.8u
m19977 VDDREF 3147 3372 VDDREF pch l=0.04u w=0.8u
m19978 VDDREF 3404 30961 VDDREF pch l=0.04u w=0.12u
m19979 VDDREF 3405 30962 VDDREF pch l=0.04u w=0.12u
m19980 VDDREF 3149 3373 VDDREF pch l=0.04u w=0.8u
m19981 3388 3295 3370 VDDREF pch l=0.04u w=0.8u
m19982 VDDREF 3150 3374 VDDREF pch l=0.04u w=0.8u
m19983 VDDREF 3151 3375 VDDREF pch l=0.04u w=0.8u
m19984 VDDREF 3153 3376 VDDREF pch l=0.04u w=0.8u
m19985 VDDREF 3154 3377 VDDREF pch l=0.04u w=0.8u
m19986 VDDREF 3155 3378 VDDREF pch l=0.04u w=0.8u
m19987 VDDREF 3157 3379 VDDREF pch l=0.04u w=0.8u
m19988 VDDREF 3158 3380 VDDREF pch l=0.04u w=0.8u
m19989 VDDREF 3317 3365 VDDREF pch l=0.04u w=0.8u
m19990 3394 3013 3381 VDDREF pch l=0.04u w=0.8u
m19991 30977 4251 3387 VDDREF pch l=0.04u w=0.12u
m19992 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m19993 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m19994 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m19995 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m19996 VDDREF 3406 30969 VDDREF pch l=0.04u w=0.12u
m19997 3395 3296 3383 VDDREF pch l=0.04u w=0.8u
m19998 3396 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m19999 3397 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20000 3398 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20001 3399 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20002 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m20003 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m20004 VDDREF 3410 30972 VDDREF pch l=0.04u w=0.12u
m20005 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m20006 3401 3360 VDDREF VDDREF pch l=0.04u w=0.8u
m20007 3402 3366 VDDREF VDDREF pch l=0.04u w=0.8u
m20008 3403 3367 VDDREF VDDREF pch l=0.04u w=0.8u
m20009 VDDREF 3203 3389 VDDREF pch l=0.04u w=0.8u
m20010 VDDREF 3208 3390 VDDREF pch l=0.04u w=0.8u
m20011 3404 3368 VDDREF VDDREF pch l=0.04u w=0.8u
m20012 3405 3369 VDDREF VDDREF pch l=0.04u w=0.8u
m20013 VDDREF 3204 3391 VDDREF pch l=0.04u w=0.8u
m20014 30980 4328 3388 VDDREF pch l=0.04u w=0.12u
m20015 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m20016 VDDREF 2854 3392 VDDREF pch l=0.04u w=0.8u
m20017 VDDREF 2856 3393 VDDREF pch l=0.04u w=0.8u
m20018 VDDREF 3386 3394 VDDREF pch l=0.04u w=0.8u
m20019 VDDREF 3070 30977 VDDREF pch l=0.04u w=0.12u
m20020 3406 3382 VDDREF VDDREF pch l=0.04u w=0.8u
m20021 30985 4328 3395 VDDREF pch l=0.04u w=0.12u
m20022 VDDREF 3434 3400 VDDREF pch l=0.04u w=0.8u
m20023 VDDREF 3432 VDDREF VDDREF pch l=0.26u w=1u
m20024 3410 3384 VDDREF VDDREF pch l=0.04u w=0.8u
m20025 3411 3288 VDDREF VDDREF pch l=0.04u w=0.8u
m20026 VDDREF 3256 3401 VDDREF pch l=0.04u w=0.8u
m20027 VDDREF 3440 30980 VDDREF pch l=0.04u w=0.12u
m20028 3413 3371 VDDREF VDDREF pch l=0.04u w=0.8u
m20029 3415 3372 VDDREF VDDREF pch l=0.04u w=0.8u
m20030 3417 3373 VDDREF VDDREF pch l=0.04u w=0.8u
m20031 3418 3374 VDDREF VDDREF pch l=0.04u w=0.8u
m20032 3419 3375 VDDREF VDDREF pch l=0.04u w=0.8u
m20033 3421 3376 VDDREF VDDREF pch l=0.04u w=0.8u
m20034 3422 3377 VDDREF VDDREF pch l=0.04u w=0.8u
m20035 3423 3378 VDDREF VDDREF pch l=0.04u w=0.8u
m20036 3425 3379 VDDREF VDDREF pch l=0.04u w=0.8u
m20037 3426 3380 VDDREF VDDREF pch l=0.04u w=0.8u
m20038 3070 3387 VDDREF VDDREF pch l=0.04u w=0.8u
m20039 3427 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m20040 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m20041 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m20042 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m20043 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m20044 VDDREF 3442 30985 VDDREF pch l=0.04u w=0.12u
m20045 3428 4328 3407 VDDREF pch l=0.04u w=0.8u
m20046 3429 4328 3408 VDDREF pch l=0.04u w=0.8u
m20047 3430 4328 3409 VDDREF pch l=0.04u w=0.8u
m20048 3431 4328 3341 VDDREF pch l=0.04u w=0.8u
m20049 3433 3433 VDDREF VDDREF pch l=0.04u w=1u
m20050 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m20051 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m20052 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m20053 VDDREF 3446 VDDREF VDDREF pch l=0.26u w=1u
m20054 3440 3388 VDDREF VDDREF pch l=0.04u w=0.8u
m20055 3436 3354 3402 VDDREF pch l=0.04u w=0.8u
m20056 3437 3355 3403 VDDREF pch l=0.04u w=0.8u
m20057 3412 3203 VDDREF VDDREF pch l=0.04u w=0.8u
m20058 VDDREF 3274 3413 VDDREF pch l=0.04u w=0.8u
m20059 3414 3208 VDDREF VDDREF pch l=0.04u w=0.8u
m20060 VDDREF 3275 3415 VDDREF pch l=0.04u w=0.8u
m20061 3438 3356 3404 VDDREF pch l=0.04u w=0.8u
m20062 3439 3357 3405 VDDREF pch l=0.04u w=0.8u
m20063 3416 3204 VDDREF VDDREF pch l=0.04u w=0.8u
m20064 VDDREF 3278 3417 VDDREF pch l=0.04u w=0.8u
m20065 VDDREF 3279 3418 VDDREF pch l=0.04u w=0.8u
m20066 VDDREF 3280 3419 VDDREF pch l=0.04u w=0.8u
m20067 3420 2854 VDDREF VDDREF pch l=0.04u w=0.8u
m20068 VDDREF 3281 3421 VDDREF pch l=0.04u w=0.8u
m20069 VDDREF 3282 3422 VDDREF pch l=0.04u w=0.8u
m20070 VDDREF 3283 3423 VDDREF pch l=0.04u w=0.8u
m20071 3424 2856 VDDREF VDDREF pch l=0.04u w=0.8u
m20072 VDDREF 3284 3425 VDDREF pch l=0.04u w=0.8u
m20073 VDDREF 3285 3426 VDDREF pch l=0.04u w=0.8u
m20074 3386 3953 VDDREF VDDREF pch l=0.04u w=0.8u
m20075 3442 3395 VDDREF VDDREF pch l=0.04u w=0.8u
m20076 3441 3358 3406 VDDREF pch l=0.04u w=0.8u
m20077 31000 3396 3428 VDDREF pch l=0.04u w=0.12u
m20078 31001 3397 3429 VDDREF pch l=0.04u w=0.12u
m20079 31002 3398 3430 VDDREF pch l=0.04u w=0.12u
m20080 31003 3399 3431 VDDREF pch l=0.04u w=0.12u
m20081 VDDREF 3484 3434 VDDREF pch l=0.04u w=0.8u
m20082 3445 3445 VDDREF VDDREF pch l=0.04u w=1u
m20083 3447 3359 3410 VDDREF pch l=0.04u w=0.8u
m20084 3435 3115 3288 VDDREF pch l=0.04u w=0.8u
m20085 3448 3302 VDDREF VDDREF pch l=0.04u w=0.8u
m20086 31006 4328 3436 VDDREF pch l=0.04u w=0.12u
m20087 31007 4328 3437 VDDREF pch l=0.04u w=0.12u
m20088 VDDREF 3204 3412 VDDREF pch l=0.04u w=0.8u
m20089 VDDREF 2024 3414 VDDREF pch l=0.04u w=0.8u
m20090 31008 4328 3438 VDDREF pch l=0.04u w=0.12u
m20091 31009 4328 3439 VDDREF pch l=0.04u w=0.12u
m20092 VDDREF FRAC[14] 3416 VDDREF pch l=0.04u w=0.8u
m20093 VDDREF 2744 3420 VDDREF pch l=0.04u w=0.8u
m20094 VDDREF FRAC[14] 3424 VDDREF pch l=0.04u w=0.8u
m20095 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m20096 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m20097 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m20098 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m20099 VDDREF 3484 3386 VDDREF pch l=0.04u w=0.8u
m20100 3450 3070 VDDREF VDDREF pch l=0.04u w=0.8u
m20101 3449 4251 3365 VDDREF pch l=0.04u w=0.8u
m20102 31014 4328 3441 VDDREF pch l=0.04u w=0.12u
m20103 VDDREF 3470 31000 VDDREF pch l=0.04u w=0.12u
m20104 VDDREF 3471 31001 VDDREF pch l=0.04u w=0.12u
m20105 VDDREF 3472 31002 VDDREF pch l=0.04u w=0.12u
m20106 VDDREF 3473 31003 VDDREF pch l=0.04u w=0.12u
m20107 VDDREF 3474 VDDREF VDDREF pch l=0.26u w=1u
m20108 VDDREF 3477 VDDREF VDDREF pch l=0.26u w=1u
m20109 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m20110 3434 4351 VDDREF VDDREF pch l=0.04u w=0.8u
m20111 VDDREF 3443 3444 VDDREF pch l=0.04u w=1u
m20112 31016 4251 3447 VDDREF pch l=0.04u w=0.12u
m20113 3115 3288 3435 VDDREF pch l=0.04u w=0.8u
m20114 VDDREF 3478 31006 VDDREF pch l=0.04u w=0.12u
m20115 VDDREF 3336 31007 VDDREF pch l=0.04u w=0.12u
m20116 VDDREF 3479 31008 VDDREF pch l=0.04u w=0.12u
m20117 VDDREF 3338 31009 VDDREF pch l=0.04u w=0.12u
m20118 3456 3321 VDDREF VDDREF pch l=0.04u w=0.8u
m20119 3458 3323 VDDREF VDDREF pch l=0.04u w=0.8u
m20120 3460 3325 VDDREF VDDREF pch l=0.04u w=0.8u
m20121 3461 3327 VDDREF VDDREF pch l=0.04u w=0.8u
m20122 3462 3328 VDDREF VDDREF pch l=0.04u w=0.8u
m20123 3464 3330 VDDREF VDDREF pch l=0.04u w=0.8u
m20124 3465 3331 VDDREF VDDREF pch l=0.04u w=0.8u
m20125 3466 3332 VDDREF VDDREF pch l=0.04u w=0.8u
m20126 3468 3334 VDDREF VDDREF pch l=0.04u w=0.8u
m20127 3469 3335 VDDREF VDDREF pch l=0.04u w=0.8u
m20128 VDDREF 3070 3450 VDDREF pch l=0.04u w=0.8u
m20129 31022 3427 3449 VDDREF pch l=0.04u w=0.12u
m20130 VDDREF 3485 31014 VDDREF pch l=0.04u w=0.12u
m20131 VDDREF 3442 3451 VDDREF pch l=0.04u w=0.8u
m20132 3470 3428 VDDREF VDDREF pch l=0.04u w=0.8u
m20133 3471 3429 VDDREF VDDREF pch l=0.04u w=0.8u
m20134 3472 3430 VDDREF VDDREF pch l=0.04u w=0.8u
m20135 3473 3431 VDDREF VDDREF pch l=0.04u w=0.8u
m20136 3475 3475 VDDREF VDDREF pch l=0.04u w=1u
m20137 3476 3476 VDDREF VDDREF pch l=0.04u w=1u
m20138 VDDREF 3490 3434 VDDREF pch l=0.04u w=0.8u
m20139 VDDREF 3453 3452 VDDREF pch l=0.04u w=1u
m20140 VDDREF 3122 31016 VDDREF pch l=0.04u w=0.12u
m20141 3478 3436 VDDREF VDDREF pch l=0.04u w=0.8u
m20142 3336 3437 VDDREF VDDREF pch l=0.04u w=0.8u
m20143 VDDREF 3491 VDDREF VDDREF pch l=0.26u w=1u
m20144 VDDREF 3494 VDDREF VDDREF pch l=0.26u w=1u
m20145 3479 3438 VDDREF VDDREF pch l=0.04u w=0.8u
m20146 3338 3439 VDDREF VDDREF pch l=0.04u w=0.8u
m20147 VDDREF 3495 VDDREF VDDREF pch l=0.26u w=1u
m20148 VDDREF 3498 VDDREF VDDREF pch l=0.26u w=1u
m20149 31025 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m20150 3454 3136 3302 VDDREF pch l=0.04u w=0.8u
m20151 3362 3500 3455 VDDREF pch l=0.04u w=0.8u
m20152 3481 3501 3457 VDDREF pch l=0.04u w=0.8u
m20153 3483 3502 3459 VDDREF pch l=0.04u w=0.8u
m20154 3086 3503 3463 VDDREF pch l=0.04u w=0.8u
m20155 3087 3504 3467 VDDREF pch l=0.04u w=0.8u
m20156 VDDREF 3505 31022 VDDREF pch l=0.04u w=0.12u
m20157 3484 3518 VDDREF VDDREF pch l=0.04u w=0.8u
m20158 3485 3441 VDDREF VDDREF pch l=0.04u w=0.8u
m20159 1321 3451 VDDREF VDDREF pch l=0.04u w=0.8u
m20160 VDDREF 3512 VDDREF VDDREF pch l=0.26u w=1u
m20161 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20162 3122 3447 VDDREF VDDREF pch l=0.04u w=0.8u
m20163 3492 3492 VDDREF VDDREF pch l=0.04u w=1u
m20164 3493 3493 VDDREF VDDREF pch l=0.04u w=1u
m20165 3496 3496 VDDREF VDDREF pch l=0.04u w=1u
m20166 3497 3497 VDDREF VDDREF pch l=0.04u w=1u
m20167 3480 3435 31025 VDDREF pch l=0.04u w=0.8u
m20168 3499 3385 VDDREF VDDREF pch l=0.04u w=0.8u
m20169 3136 3302 3454 VDDREF pch l=0.04u w=0.8u
m20170 3500 3455 3362 VDDREF pch l=0.04u w=0.8u
m20171 3501 3457 3481 VDDREF pch l=0.04u w=0.8u
m20172 3502 3459 3483 VDDREF pch l=0.04u w=0.8u
m20173 3503 3463 3086 VDDREF pch l=0.04u w=0.8u
m20174 3504 3467 3087 VDDREF pch l=0.04u w=0.8u
m20175 3363 3145 3321 VDDREF pch l=0.04u w=0.8u
m20176 3482 3147 3323 VDDREF pch l=0.04u w=0.8u
m20177 3337 3149 3325 VDDREF pch l=0.04u w=0.8u
m20178 3315 3150 3327 VDDREF pch l=0.04u w=0.8u
m20179 3408 3151 3328 VDDREF pch l=0.04u w=0.8u
m20180 3253 3153 3330 VDDREF pch l=0.04u w=0.8u
m20181 3352 3154 3331 VDDREF pch l=0.04u w=0.8u
m20182 3341 3155 3332 VDDREF pch l=0.04u w=0.8u
m20183 3254 3157 3334 VDDREF pch l=0.04u w=0.8u
m20184 3353 3158 3335 VDDREF pch l=0.04u w=0.8u
m20185 3505 3449 VDDREF VDDREF pch l=0.04u w=0.8u
m20186 VDDREF 3518 3484 VDDREF pch l=0.04u w=0.8u
m20187 3506 3450 VDDREF VDDREF pch l=0.04u w=0.8u
m20188 3511 3511 VDDREF VDDREF pch l=0.04u w=1u
m20189 3507 3396 3470 VDDREF pch l=0.04u w=0.8u
m20190 3508 3397 3471 VDDREF pch l=0.04u w=0.8u
m20191 3509 3398 3472 VDDREF pch l=0.04u w=0.8u
m20192 3510 3399 3473 VDDREF pch l=0.04u w=0.8u
m20193 VDDREF 3486 3487 VDDREF pch l=0.04u w=1u
m20194 VDDREF 3489 3488 VDDREF pch l=0.04u w=1u
m20195 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20196 VDDREF 3523 3490 VDDREF pch l=0.04u w=0.8u
m20197 3145 3321 3363 VDDREF pch l=0.04u w=0.8u
m20198 3147 3323 3482 VDDREF pch l=0.04u w=0.8u
m20199 3149 3325 3337 VDDREF pch l=0.04u w=0.8u
m20200 3150 3327 3315 VDDREF pch l=0.04u w=0.8u
m20201 3151 3328 3408 VDDREF pch l=0.04u w=0.8u
m20202 3153 3330 3253 VDDREF pch l=0.04u w=0.8u
m20203 3154 3331 3352 VDDREF pch l=0.04u w=0.8u
m20204 3155 3332 3341 VDDREF pch l=0.04u w=0.8u
m20205 3157 3334 3254 VDDREF pch l=0.04u w=0.8u
m20206 3158 3335 3353 VDDREF pch l=0.04u w=0.8u
m20207 VDDREF 2969 3506 VDDREF pch l=0.04u w=0.8u
m20208 3519 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20209 3520 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20210 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20211 31053 4328 3507 VDDREF pch l=0.04u w=0.12u
m20212 31054 4328 3508 VDDREF pch l=0.04u w=0.12u
m20213 31055 4328 3509 VDDREF pch l=0.04u w=0.12u
m20214 31056 4328 3510 VDDREF pch l=0.04u w=0.12u
m20215 3524 3122 VDDREF VDDREF pch l=0.04u w=0.8u
m20216 3525 2491 VDDREF VDDREF pch l=0.04u w=0.8u
m20217 3526 110 VDDREF VDDREF pch l=0.04u w=0.8u
m20218 VDDREF 3500 3513 VDDREF pch l=0.04u w=0.8u
m20219 VDDREF 3501 3514 VDDREF pch l=0.04u w=0.8u
m20220 VDDREF 3502 3515 VDDREF pch l=0.04u w=0.8u
m20221 VDDREF 3503 3516 VDDREF pch l=0.04u w=0.8u
m20222 VDDREF 3504 3517 VDDREF pch l=0.04u w=0.8u
m20223 3506 3484 VDDREF VDDREF pch l=0.04u w=0.8u
m20224 3527 3427 3505 VDDREF pch l=0.04u w=0.8u
m20225 VDDREF 3556 3518 VDDREF pch l=0.04u w=0.8u
m20226 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20227 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20228 VDDREF 3553 31053 VDDREF pch l=0.04u w=0.12u
m20229 VDDREF 3339 31054 VDDREF pch l=0.04u w=0.12u
m20230 VDDREF 3554 31055 VDDREF pch l=0.04u w=0.12u
m20231 VDDREF 3342 31056 VDDREF pch l=0.04u w=0.12u
m20232 VDDREF 3522 3521 VDDREF pch l=0.04u w=1u
m20233 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20234 3523 4064 VDDREF VDDREF pch l=0.04u w=0.8u
m20235 VDDREF 3122 3524 VDDREF pch l=0.04u w=0.8u
m20236 VDDREF 2739 3525 VDDREF pch l=0.04u w=0.8u
m20237 VDDREF 1023 3526 VDDREF pch l=0.04u w=0.8u
m20238 VDDREF 3528 3529 VDDREF pch l=0.04u w=1u
m20239 VDDREF 3531 3530 VDDREF pch l=0.04u w=1u
m20240 3539 3610 VDDREF VDDREF pch l=0.04u w=0.8u
m20241 3540 1935 VDDREF VDDREF pch l=0.04u w=0.8u
m20242 3541 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m20243 3542 2616 VDDREF VDDREF pch l=0.04u w=0.8u
m20244 VDDREF 3532 3533 VDDREF pch l=0.04u w=1u
m20245 VDDREF 3535 3534 VDDREF pch l=0.04u w=1u
m20246 3543 FRAC[11] VDDREF VDDREF pch l=0.04u w=0.8u
m20247 VDDREF 3582 3536 VDDREF pch l=0.04u w=0.8u
m20248 3544 3611 VDDREF VDDREF pch l=0.04u w=0.8u
m20249 3545 3622 VDDREF VDDREF pch l=0.04u w=0.8u
m20250 3546 3588 VDDREF VDDREF pch l=0.04u w=0.8u
m20251 3547 3536 VDDREF VDDREF pch l=0.04u w=0.8u
m20252 3548 3623 VDDREF VDDREF pch l=0.04u w=0.8u
m20253 3549 FRAC[11] VDDREF VDDREF pch l=0.04u w=0.8u
m20254 3550 3536 VDDREF VDDREF pch l=0.04u w=0.8u
m20255 31071 4251 3527 VDDREF pch l=0.04u w=0.12u
m20256 31072 3518 VDDREF VDDREF pch l=0.04u w=0.12u
m20257 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20258 VDDREF 3538 3537 VDDREF pch l=0.04u w=1u
m20259 3551 4328 3485 VDDREF pch l=0.04u w=0.8u
m20260 3552 4328 3442 VDDREF pch l=0.04u w=0.8u
m20261 3553 3507 VDDREF VDDREF pch l=0.04u w=0.8u
m20262 3339 3508 VDDREF VDDREF pch l=0.04u w=0.8u
m20263 3554 3509 VDDREF VDDREF pch l=0.04u w=0.8u
m20264 3342 3510 VDDREF VDDREF pch l=0.04u w=0.8u
m20265 VDDREF 3565 3523 VDDREF pch l=0.04u w=0.8u
m20266 3525 3016 VDDREF VDDREF pch l=0.04u w=0.8u
m20267 3183 3693 VDDREF VDDREF pch l=0.04u w=0.8u
m20268 VDDREF 3608 3539 VDDREF pch l=0.04u w=0.8u
m20269 3185 3695 VDDREF VDDREF pch l=0.04u w=0.8u
m20270 VDDREF 3609 3540 VDDREF pch l=0.04u w=0.8u
m20271 VDDREF 3761 3541 VDDREF pch l=0.04u w=0.8u
m20272 VDDREF 3762 3542 VDDREF pch l=0.04u w=0.8u
m20273 3187 3697 VDDREF VDDREF pch l=0.04u w=0.8u
m20274 VDDREF 3610 3543 VDDREF pch l=0.04u w=0.8u
m20275 VDDREF 131 3544 VDDREF pch l=0.04u w=0.8u
m20276 VDDREF 3611 3545 VDDREF pch l=0.04u w=0.8u
m20277 3191 3701 VDDREF VDDREF pch l=0.04u w=0.8u
m20278 VDDREF 3612 3546 VDDREF pch l=0.04u w=0.8u
m20279 VDDREF 3589 3547 VDDREF pch l=0.04u w=0.8u
m20280 VDDREF 3613 3548 VDDREF pch l=0.04u w=0.8u
m20281 3195 3705 VDDREF VDDREF pch l=0.04u w=0.8u
m20282 VDDREF 3614 3549 VDDREF pch l=0.04u w=0.8u
m20283 VDDREF FBDIV[11] 3550 VDDREF pch l=0.04u w=0.8u
m20284 VDDREF 3199 31071 VDDREF pch l=0.04u w=0.12u
m20285 3556 4251 31072 VDDREF pch l=0.04u w=0.12u
m20286 3555 3506 VDDREF VDDREF pch l=0.04u w=0.8u
m20287 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20288 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20289 VDDREF 3679 VDDREF VDDREF pch l=0.26u w=1u
m20290 31083 3519 3551 VDDREF pch l=0.04u w=0.12u
m20291 31084 3520 3552 VDDREF pch l=0.04u w=0.12u
m20292 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20293 3557 3567 VDDREF VDDREF pch l=0.04u w=0.8u
m20294 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20295 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20296 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20297 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20298 3558 1023 VDDREF VDDREF pch l=0.04u w=0.8u
m20299 VDDREF 3591 3183 VDDREF pch l=0.04u w=0.8u
m20300 VDDREF 3593 3185 VDDREF pch l=0.04u w=0.8u
m20301 VDDREF 3595 3187 VDDREF pch l=0.04u w=0.8u
m20302 VDDREF 3600 3191 VDDREF pch l=0.04u w=0.8u
m20303 VDDREF 3604 3195 VDDREF pch l=0.04u w=0.8u
m20304 3199 3527 VDDREF VDDREF pch l=0.04u w=0.8u
m20305 3559 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20306 3560 3660 3556 VDDREF pch l=0.04u w=0.8u
m20307 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20308 VDDREF 3690 VDDREF VDDREF pch l=0.26u w=1u
m20309 VDDREF 3584 31083 VDDREF pch l=0.04u w=0.12u
m20310 VDDREF 3585 31084 VDDREF pch l=0.04u w=0.12u
m20311 3561 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20312 3562 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20313 3563 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20314 3564 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20315 3565 3619 VDDREF VDDREF pch l=0.04u w=0.8u
m20316 3566 3590 3557 VDDREF pch l=0.04u w=0.8u
m20317 3568 3525 VDDREF VDDREF pch l=0.04u w=0.8u
m20318 3570 3608 VDDREF VDDREF pch l=0.04u w=0.8u
m20319 3571 3609 VDDREF VDDREF pch l=0.04u w=0.8u
m20320 3572 3541 VDDREF VDDREF pch l=0.04u w=0.8u
m20321 3573 3542 VDDREF VDDREF pch l=0.04u w=0.8u
m20322 3574 3610 VDDREF VDDREF pch l=0.04u w=0.8u
m20323 3575 131 VDDREF VDDREF pch l=0.04u w=0.8u
m20324 3576 3611 VDDREF VDDREF pch l=0.04u w=0.8u
m20325 3577 3612 VDDREF VDDREF pch l=0.04u w=0.8u
m20326 3578 3589 VDDREF VDDREF pch l=0.04u w=0.8u
m20327 3579 3613 VDDREF VDDREF pch l=0.04u w=0.8u
m20328 3580 3614 VDDREF VDDREF pch l=0.04u w=0.8u
m20329 3581 FBDIV[11] VDDREF VDDREF pch l=0.04u w=0.8u
m20330 3583 3555 VDDREF VDDREF pch l=0.04u w=0.8u
m20331 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20332 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20333 VDDREF 3679 VDDREF VDDREF pch l=0.26u w=1u
m20334 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20335 3584 3551 VDDREF VDDREF pch l=0.04u w=0.8u
m20336 3585 3552 VDDREF VDDREF pch l=0.04u w=0.8u
m20337 VDDREF 3619 3565 VDDREF pch l=0.04u w=0.8u
m20338 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20339 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20340 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20341 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20342 3590 3557 3566 VDDREF pch l=0.04u w=0.8u
m20343 3569 110 1023 VDDREF pch l=0.04u w=0.8u
m20344 3591 3455 VDDREF VDDREF pch l=0.04u w=0.8u
m20345 3593 3457 VDDREF VDDREF pch l=0.04u w=0.8u
m20346 3595 3459 VDDREF VDDREF pch l=0.04u w=0.8u
m20347 3600 3463 VDDREF VDDREF pch l=0.04u w=0.8u
m20348 3604 3467 VDDREF VDDREF pch l=0.04u w=0.8u
m20349 3607 3199 VDDREF VDDREF pch l=0.04u w=0.8u
m20350 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20351 VDDREF 3690 VDDREF VDDREF pch l=0.26u w=1u
m20352 3597 4328 3582 VDDREF pch l=0.04u w=0.8u
m20353 VDDREF 3634 3560 VDDREF pch l=0.04u w=0.8u
m20354 VDDREF 3953 3583 VDDREF pch l=0.04u w=0.8u
m20355 3615 4328 3586 VDDREF pch l=0.04u w=0.8u
m20356 3616 4328 3587 VDDREF pch l=0.04u w=0.8u
m20357 3617 4328 3588 VDDREF pch l=0.04u w=0.8u
m20358 3618 4328 3589 VDDREF pch l=0.04u w=0.8u
m20359 3620 3568 VDDREF VDDREF pch l=0.04u w=0.8u
m20360 110 1023 3569 VDDREF pch l=0.04u w=0.8u
m20361 VDDREF 3500 3591 VDDREF pch l=0.04u w=0.8u
m20362 VDDREF 3501 3593 VDDREF pch l=0.04u w=0.8u
m20363 VDDREF 3502 3595 VDDREF pch l=0.04u w=0.8u
m20364 VDDREF 3503 3600 VDDREF pch l=0.04u w=0.8u
m20365 VDDREF 3504 3604 VDDREF pch l=0.04u w=0.8u
m20366 VDDREF 3199 3607 VDDREF pch l=0.04u w=0.8u
m20367 3624 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20368 3625 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20369 3592 3610 3608 VDDREF pch l=0.04u w=0.8u
m20370 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20371 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20372 3594 1935 3609 VDDREF pch l=0.04u w=0.8u
m20373 3626 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20374 3627 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20375 3596 FRAC[11] 3610 VDDREF pch l=0.04u w=0.8u
m20376 31140 3559 3597 VDDREF pch l=0.04u w=0.12u
m20377 3598 3611 131 VDDREF pch l=0.04u w=0.8u
m20378 3599 3622 3611 VDDREF pch l=0.04u w=0.8u
m20379 3601 3588 3612 VDDREF pch l=0.04u w=0.8u
m20380 3602 3536 3589 VDDREF pch l=0.04u w=0.8u
m20381 3603 3623 3613 VDDREF pch l=0.04u w=0.8u
m20382 3605 FRAC[11] 3614 VDDREF pch l=0.04u w=0.8u
m20383 3606 3536 FBDIV[11] VDDREF pch l=0.04u w=0.8u
m20384 31143 3560 VDDREF VDDREF pch l=0.04u w=0.12u
m20385 VDDREF 3679 VDDREF VDDREF pch l=0.26u w=1u
m20386 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20387 3628 3519 3584 VDDREF pch l=0.04u w=0.8u
m20388 3629 3520 3585 VDDREF pch l=0.04u w=0.8u
m20389 31294 3561 3615 VDDREF pch l=0.04u w=0.12u
m20390 31295 3562 3616 VDDREF pch l=0.04u w=0.12u
m20391 31296 3563 3617 VDDREF pch l=0.04u w=0.12u
m20392 31297 3564 3618 VDDREF pch l=0.04u w=0.12u
m20393 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20394 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20395 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20396 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20397 VDDREF 3659 3619 VDDREF pch l=0.04u w=0.8u
m20398 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20399 VDDREF 3690 VDDREF VDDREF pch l=0.26u w=1u
m20400 VDDREF 3288 3620 VDDREF pch l=0.04u w=0.8u
m20401 3610 3608 3592 VDDREF pch l=0.04u w=0.8u
m20402 1935 3609 3594 VDDREF pch l=0.04u w=0.8u
m20403 FRAC[11] 3610 3596 VDDREF pch l=0.04u w=0.8u
m20404 VDDREF 3641 31140 VDDREF pch l=0.04u w=0.12u
m20405 3611 131 3598 VDDREF pch l=0.04u w=0.8u
m20406 3622 3611 3599 VDDREF pch l=0.04u w=0.8u
m20407 3588 3612 3601 VDDREF pch l=0.04u w=0.8u
m20408 3536 3589 3602 VDDREF pch l=0.04u w=0.8u
m20409 3623 3613 3603 VDDREF pch l=0.04u w=0.8u
m20410 FRAC[11] 3614 3605 VDDREF pch l=0.04u w=0.8u
m20411 3536 FBDIV[11] 3606 VDDREF pch l=0.04u w=0.8u
m20412 3634 3660 31143 VDDREF pch l=0.04u w=0.12u
m20413 3635 3583 VDDREF VDDREF pch l=0.04u w=0.8u
m20414 31305 4328 3628 VDDREF pch l=0.04u w=0.12u
m20415 31306 4328 3629 VDDREF pch l=0.04u w=0.12u
m20416 VDDREF 3655 31294 VDDREF pch l=0.04u w=0.12u
m20417 VDDREF 3656 31295 VDDREF pch l=0.04u w=0.12u
m20418 VDDREF 3657 31296 VDDREF pch l=0.04u w=0.12u
m20419 VDDREF 3658 31297 VDDREF pch l=0.04u w=0.12u
m20420 31462 3619 VDDREF VDDREF pch l=0.04u w=0.12u
m20421 3636 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m20422 3620 2630 VDDREF VDDREF pch l=0.04u w=0.8u
m20423 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20424 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20425 VDDREF 3679 VDDREF VDDREF pch l=0.26u w=1u
m20426 3630 3569 VDDREF VDDREF pch l=0.04u w=0.8u
m20427 3500 3478 3479 VDDREF pch l=0.04u w=0.8u
m20428 3501 3483 1998 VDDREF pch l=0.04u w=0.8u
m20429 3502 3479 FRAC[13] VDDREF pch l=0.04u w=0.8u
m20430 3641 3597 VDDREF VDDREF pch l=0.04u w=0.8u
m20431 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20432 3503 3201 3087 VDDREF pch l=0.04u w=0.8u
m20433 3504 3202 FRAC[13] VDDREF pch l=0.04u w=0.8u
m20434 3642 4251 3634 VDDREF pch l=0.04u w=0.8u
m20435 3643 3484 VDDREF VDDREF pch l=0.04u w=0.8u
m20436 3637 4328 3632 VDDREF pch l=0.04u w=0.8u
m20437 3638 4328 3633 VDDREF pch l=0.04u w=0.8u
m20438 3639 4328 3572 VDDREF pch l=0.04u w=0.8u
m20439 3640 4328 3573 VDDREF pch l=0.04u w=0.8u
m20440 3654 3661 3635 VDDREF pch l=0.04u w=0.8u
m20441 VDDREF 3662 31305 VDDREF pch l=0.04u w=0.12u
m20442 VDDREF 3663 31306 VDDREF pch l=0.04u w=0.12u
m20443 3655 3615 VDDREF VDDREF pch l=0.04u w=0.8u
m20444 3656 3616 VDDREF VDDREF pch l=0.04u w=0.8u
m20445 3657 3617 VDDREF VDDREF pch l=0.04u w=0.8u
m20446 3658 3618 VDDREF VDDREF pch l=0.04u w=0.8u
m20447 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20448 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20449 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20450 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20451 3659 4251 31462 VDDREF pch l=0.04u w=0.12u
m20452 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20453 VDDREF 3690 VDDREF VDDREF pch l=0.26u w=1u
m20454 VDDREF 3401 3630 VDDREF pch l=0.04u w=0.8u
m20455 3478 3479 3500 VDDREF pch l=0.04u w=0.8u
m20456 3483 1998 3501 VDDREF pch l=0.04u w=0.8u
m20457 3479 FRAC[13] 3502 VDDREF pch l=0.04u w=0.8u
m20458 3201 3087 3503 VDDREF pch l=0.04u w=0.8u
m20459 3202 FRAC[13] 3504 VDDREF pch l=0.04u w=0.8u
m20460 31468 3624 3637 VDDREF pch l=0.04u w=0.12u
m20461 31469 3625 3638 VDDREF pch l=0.04u w=0.12u
m20462 3644 3592 VDDREF VDDREF pch l=0.04u w=0.8u
m20463 3645 3594 VDDREF VDDREF pch l=0.04u w=0.8u
m20464 31470 3626 3639 VDDREF pch l=0.04u w=0.12u
m20465 31471 3627 3640 VDDREF pch l=0.04u w=0.12u
m20466 3646 3596 VDDREF VDDREF pch l=0.04u w=0.8u
m20467 3647 3598 VDDREF VDDREF pch l=0.04u w=0.8u
m20468 3648 3599 VDDREF VDDREF pch l=0.04u w=0.8u
m20469 3649 3601 VDDREF VDDREF pch l=0.04u w=0.8u
m20470 3650 3602 VDDREF VDDREF pch l=0.04u w=0.8u
m20471 3651 3603 VDDREF VDDREF pch l=0.04u w=0.8u
m20472 3652 3605 VDDREF VDDREF pch l=0.04u w=0.8u
m20473 3653 3606 VDDREF VDDREF pch l=0.04u w=0.8u
m20474 3661 3635 3654 VDDREF pch l=0.04u w=0.8u
m20475 3662 3628 VDDREF VDDREF pch l=0.04u w=0.8u
m20476 3663 3629 VDDREF VDDREF pch l=0.04u w=0.8u
m20477 3664 3756 3659 VDDREF pch l=0.04u w=0.8u
m20478 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20479 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20480 VDDREF 3679 VDDREF VDDREF pch l=0.26u w=1u
m20481 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20482 3665 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m20483 3666 3499 VDDREF VDDREF pch l=0.04u w=0.8u
m20484 VDDREF 3681 31468 VDDREF pch l=0.04u w=0.12u
m20485 VDDREF 3682 31469 VDDREF pch l=0.04u w=0.12u
m20486 VDDREF 3413 3644 VDDREF pch l=0.04u w=0.8u
m20487 VDDREF 3415 3645 VDDREF pch l=0.04u w=0.8u
m20488 VDDREF 3683 31470 VDDREF pch l=0.04u w=0.12u
m20489 VDDREF 3684 31471 VDDREF pch l=0.04u w=0.12u
m20490 VDDREF 3417 3646 VDDREF pch l=0.04u w=0.8u
m20491 3667 3559 3641 VDDREF pch l=0.04u w=0.8u
m20492 VDDREF 3418 3647 VDDREF pch l=0.04u w=0.8u
m20493 VDDREF 3419 3648 VDDREF pch l=0.04u w=0.8u
m20494 VDDREF 3421 3649 VDDREF pch l=0.04u w=0.8u
m20495 VDDREF 3422 3650 VDDREF pch l=0.04u w=0.8u
m20496 VDDREF 3423 3651 VDDREF pch l=0.04u w=0.8u
m20497 VDDREF 3425 3652 VDDREF pch l=0.04u w=0.8u
m20498 VDDREF 3426 3653 VDDREF pch l=0.04u w=0.8u
m20499 VDDREF 4251 3660 VDDREF pch l=0.04u w=0.8u
m20500 3673 3607 VDDREF VDDREF pch l=0.04u w=0.8u
m20501 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20502 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20503 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20504 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20505 3674 3561 3655 VDDREF pch l=0.04u w=0.8u
m20506 3675 3562 3656 VDDREF pch l=0.04u w=0.8u
m20507 3676 3563 3657 VDDREF pch l=0.04u w=0.8u
m20508 3677 3564 3658 VDDREF pch l=0.04u w=0.8u
m20509 VDDREF 3687 VDDREF VDDREF pch l=0.26u w=1u
m20510 VDDREF 3690 VDDREF VDDREF pch l=0.26u w=1u
m20511 3678 3678 VDDREF VDDREF pch l=0.04u w=1u
m20512 VDDREF 616 3665 VDDREF pch l=0.04u w=0.8u
m20513 VDDREF 3620 3666 VDDREF pch l=0.04u w=0.8u
m20514 3680 3630 VDDREF VDDREF pch l=0.04u w=0.8u
m20515 3681 3637 VDDREF VDDREF pch l=0.04u w=0.8u
m20516 3682 3638 VDDREF VDDREF pch l=0.04u w=0.8u
m20517 VDDREF 3478 3668 VDDREF pch l=0.04u w=0.8u
m20518 VDDREF 3483 3669 VDDREF pch l=0.04u w=0.8u
m20519 3683 3639 VDDREF VDDREF pch l=0.04u w=0.8u
m20520 3684 3640 VDDREF VDDREF pch l=0.04u w=0.8u
m20521 VDDREF 3479 3670 VDDREF pch l=0.04u w=0.8u
m20522 31517 4328 3667 VDDREF pch l=0.04u w=0.12u
m20523 VDDREF 3201 3671 VDDREF pch l=0.04u w=0.8u
m20524 VDDREF 3202 3672 VDDREF pch l=0.04u w=0.8u
m20525 VDDREF 3017 3673 VDDREF pch l=0.04u w=0.8u
m20526 3685 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20527 3686 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20528 31669 4328 3674 VDDREF pch l=0.04u w=0.12u
m20529 31670 4328 3675 VDDREF pch l=0.04u w=0.12u
m20530 31671 4328 3676 VDDREF pch l=0.04u w=0.12u
m20531 31672 4328 3677 VDDREF pch l=0.04u w=0.12u
m20532 3688 3688 VDDREF VDDREF pch l=0.04u w=1u
m20533 3689 3689 VDDREF VDDREF pch l=0.04u w=1u
m20534 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20535 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20536 VDDREF 3722 3664 VDDREF pch l=0.04u w=0.8u
m20537 VDDREF 3712 VDDREF VDDREF pch l=0.26u w=1u
m20538 VDDREF 3526 3680 VDDREF pch l=0.04u w=0.8u
m20539 VDDREF 3719 31517 VDDREF pch l=0.04u w=0.12u
m20540 3673 4351 VDDREF VDDREF pch l=0.04u w=0.8u
m20541 3694 3644 VDDREF VDDREF pch l=0.04u w=0.8u
m20542 3696 3645 VDDREF VDDREF pch l=0.04u w=0.8u
m20543 3698 3646 VDDREF VDDREF pch l=0.04u w=0.8u
m20544 3699 3647 VDDREF VDDREF pch l=0.04u w=0.8u
m20545 3700 3648 VDDREF VDDREF pch l=0.04u w=0.8u
m20546 3702 3649 VDDREF VDDREF pch l=0.04u w=0.8u
m20547 3703 3650 VDDREF VDDREF pch l=0.04u w=0.8u
m20548 3704 3651 VDDREF VDDREF pch l=0.04u w=0.8u
m20549 3706 3652 VDDREF VDDREF pch l=0.04u w=0.8u
m20550 3707 3653 VDDREF VDDREF pch l=0.04u w=0.8u
m20551 3642 3764 VDDREF VDDREF pch l=0.04u w=0.8u
m20552 3708 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m20553 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20554 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20555 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20556 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20557 VDDREF 3612 31669 VDDREF pch l=0.04u w=0.12u
m20558 VDDREF 3611 31670 VDDREF pch l=0.04u w=0.12u
m20559 VDDREF 3614 31671 VDDREF pch l=0.04u w=0.12u
m20560 VDDREF 3613 31672 VDDREF pch l=0.04u w=0.12u
m20561 31833 3664 VDDREF VDDREF pch l=0.04u w=0.12u
m20562 3711 3711 VDDREF VDDREF pch l=0.04u w=1u
m20563 VDDREF 3692 3691 VDDREF pch l=0.04u w=1u
m20564 3713 3636 VDDREF VDDREF pch l=0.04u w=0.8u
m20565 3714 2508 VDDREF VDDREF pch l=0.04u w=0.8u
m20566 3719 3667 VDDREF VDDREF pch l=0.04u w=0.8u
m20567 3715 3624 3681 VDDREF pch l=0.04u w=0.8u
m20568 3716 3625 3682 VDDREF pch l=0.04u w=0.8u
m20569 3693 3478 VDDREF VDDREF pch l=0.04u w=0.8u
m20570 VDDREF 3539 3694 VDDREF pch l=0.04u w=0.8u
m20571 3695 3483 VDDREF VDDREF pch l=0.04u w=0.8u
m20572 VDDREF 3540 3696 VDDREF pch l=0.04u w=0.8u
m20573 3717 3626 3683 VDDREF pch l=0.04u w=0.8u
m20574 3718 3627 3684 VDDREF pch l=0.04u w=0.8u
m20575 3697 3479 VDDREF VDDREF pch l=0.04u w=0.8u
m20576 VDDREF 3543 3698 VDDREF pch l=0.04u w=0.8u
m20577 VDDREF 3544 3699 VDDREF pch l=0.04u w=0.8u
m20578 VDDREF 3545 3700 VDDREF pch l=0.04u w=0.8u
m20579 3701 3201 VDDREF VDDREF pch l=0.04u w=0.8u
m20580 VDDREF 3546 3702 VDDREF pch l=0.04u w=0.8u
m20581 VDDREF 3547 3703 VDDREF pch l=0.04u w=0.8u
m20582 VDDREF 3548 3704 VDDREF pch l=0.04u w=0.8u
m20583 3705 3202 VDDREF VDDREF pch l=0.04u w=0.8u
m20584 VDDREF 3549 3706 VDDREF pch l=0.04u w=0.8u
m20585 VDDREF 3550 3707 VDDREF pch l=0.04u w=0.8u
m20586 VDDREF 3800 3642 VDDREF pch l=0.04u w=0.8u
m20587 3720 4328 3662 VDDREF pch l=0.04u w=0.8u
m20588 3721 4328 3663 VDDREF pch l=0.04u w=0.8u
m20589 3612 3674 VDDREF VDDREF pch l=0.04u w=0.8u
m20590 3611 3675 VDDREF VDDREF pch l=0.04u w=0.8u
m20591 3614 3676 VDDREF VDDREF pch l=0.04u w=0.8u
m20592 3613 3677 VDDREF VDDREF pch l=0.04u w=0.8u
m20593 VDDREF 3728 VDDREF VDDREF pch l=0.26u w=1u
m20594 VDDREF 3731 VDDREF VDDREF pch l=0.26u w=1u
m20595 3722 3756 31833 VDDREF pch l=0.04u w=0.12u
m20596 VDDREF 3709 3710 VDDREF pch l=0.04u w=1u
m20597 VDDREF 3566 3713 VDDREF pch l=0.04u w=0.8u
m20598 VDDREF 3180 3714 VDDREF pch l=0.04u w=0.8u
m20599 3725 3569 VDDREF VDDREF pch l=0.04u w=0.8u
m20600 31871 4328 3715 VDDREF pch l=0.04u w=0.12u
m20601 31872 4328 3716 VDDREF pch l=0.04u w=0.12u
m20602 VDDREF 3479 3693 VDDREF pch l=0.04u w=0.8u
m20603 VDDREF 1998 3695 VDDREF pch l=0.04u w=0.8u
m20604 31873 4328 3717 VDDREF pch l=0.04u w=0.12u
m20605 31874 4328 3718 VDDREF pch l=0.04u w=0.12u
m20606 VDDREF FRAC[13] 3697 VDDREF pch l=0.04u w=0.8u
m20607 VDDREF 3087 3701 VDDREF pch l=0.04u w=0.8u
m20608 VDDREF FRAC[13] 3705 VDDREF pch l=0.04u w=0.8u
m20609 3642 3800 VDDREF VDDREF pch l=0.04u w=0.8u
m20610 3726 3673 VDDREF VDDREF pch l=0.04u w=0.8u
m20611 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20612 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20613 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20614 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20615 3727 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m20616 31876 3685 3720 VDDREF pch l=0.04u w=0.12u
m20617 31877 3686 3721 VDDREF pch l=0.04u w=0.12u
m20618 3729 3729 VDDREF VDDREF pch l=0.04u w=1u
m20619 3730 3730 VDDREF VDDREF pch l=0.04u w=1u
m20620 3732 4251 3722 VDDREF pch l=0.04u w=0.8u
m20621 VDDREF 3849 VDDREF VDDREF pch l=0.26u w=1u
m20622 VDDREF 3724 3723 VDDREF pch l=0.04u w=1u
m20623 3735 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m20624 VDDREF 3759 31871 VDDREF pch l=0.04u w=0.12u
m20625 VDDREF 3608 31872 VDDREF pch l=0.04u w=0.12u
m20626 VDDREF 3760 31873 VDDREF pch l=0.04u w=0.12u
m20627 VDDREF 3610 31874 VDDREF pch l=0.04u w=0.12u
m20628 VDDREF 3764 3642 VDDREF pch l=0.04u w=0.8u
m20629 3738 3592 VDDREF VDDREF pch l=0.04u w=0.8u
m20630 3740 3594 VDDREF VDDREF pch l=0.04u w=0.8u
m20631 3742 3596 VDDREF VDDREF pch l=0.04u w=0.8u
m20632 3743 3598 VDDREF VDDREF pch l=0.04u w=0.8u
m20633 3744 3599 VDDREF VDDREF pch l=0.04u w=0.8u
m20634 3746 3601 VDDREF VDDREF pch l=0.04u w=0.8u
m20635 3747 3602 VDDREF VDDREF pch l=0.04u w=0.8u
m20636 3748 3603 VDDREF VDDREF pch l=0.04u w=0.8u
m20637 3750 3605 VDDREF VDDREF pch l=0.04u w=0.8u
m20638 3751 3606 VDDREF VDDREF pch l=0.04u w=0.8u
m20639 VDDREF 2245 3727 VDDREF pch l=0.04u w=0.8u
m20640 VDDREF 3766 31876 VDDREF pch l=0.04u w=0.12u
m20641 VDDREF 3767 31877 VDDREF pch l=0.04u w=0.12u
m20642 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20643 VDDREF 3733 3734 VDDREF pch l=0.04u w=1u
m20644 3757 3713 VDDREF VDDREF pch l=0.04u w=0.8u
m20645 VDDREF 3180 3735 VDDREF pch l=0.04u w=0.8u
m20646 3758 3180 VDDREF VDDREF pch l=0.04u w=0.8u
m20647 3759 3715 VDDREF VDDREF pch l=0.04u w=0.8u
m20648 3608 3716 VDDREF VDDREF pch l=0.04u w=0.8u
m20649 VDDREF 3769 VDDREF VDDREF pch l=0.26u w=1u
m20650 VDDREF 3772 VDDREF VDDREF pch l=0.26u w=1u
m20651 3760 3717 VDDREF VDDREF pch l=0.04u w=0.8u
m20652 3610 3718 VDDREF VDDREF pch l=0.04u w=0.8u
m20653 VDDREF 3773 VDDREF VDDREF pch l=0.26u w=1u
m20654 VDDREF 3776 VDDREF VDDREF pch l=0.26u w=1u
m20655 3736 3401 3569 VDDREF pch l=0.04u w=0.8u
m20656 3632 3777 3737 VDDREF pch l=0.04u w=0.8u
m20657 3761 3778 3739 VDDREF pch l=0.04u w=0.8u
m20658 3763 3779 3741 VDDREF pch l=0.04u w=0.8u
m20659 3407 3780 3745 VDDREF pch l=0.04u w=0.8u
m20660 3409 3781 3749 VDDREF pch l=0.04u w=0.8u
m20661 3765 3726 VDDREF VDDREF pch l=0.04u w=0.8u
m20662 3766 3720 VDDREF VDDREF pch l=0.04u w=0.8u
m20663 3767 3721 VDDREF VDDREF pch l=0.04u w=0.8u
m20664 VDDREF 3752 3753 VDDREF pch l=0.04u w=1u
m20665 VDDREF 3755 3754 VDDREF pch l=0.04u w=1u
m20666 VDDREF 3849 VDDREF VDDREF pch l=0.26u w=1u
m20667 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20668 VDDREF 4251 3756 VDDREF pch l=0.04u w=0.8u
m20669 VDDREF 3665 3757 VDDREF pch l=0.04u w=0.8u
m20670 3770 3770 VDDREF VDDREF pch l=0.04u w=1u
m20671 3771 3771 VDDREF VDDREF pch l=0.04u w=1u
m20672 3774 3774 VDDREF VDDREF pch l=0.04u w=1u
m20673 3775 3775 VDDREF VDDREF pch l=0.04u w=1u
m20674 3401 3569 3736 VDDREF pch l=0.04u w=0.8u
m20675 3777 3737 3632 VDDREF pch l=0.04u w=0.8u
m20676 3778 3739 3761 VDDREF pch l=0.04u w=0.8u
m20677 3779 3741 3763 VDDREF pch l=0.04u w=0.8u
m20678 3780 3745 3407 VDDREF pch l=0.04u w=0.8u
m20679 3781 3749 3409 VDDREF pch l=0.04u w=0.8u
m20680 3764 3862 VDDREF VDDREF pch l=0.04u w=0.8u
m20681 VDDREF 3643 3765 VDDREF pch l=0.04u w=0.8u
m20682 3633 3413 3592 VDDREF pch l=0.04u w=0.8u
m20683 3762 3415 3594 VDDREF pch l=0.04u w=0.8u
m20684 3609 3417 3596 VDDREF pch l=0.04u w=0.8u
m20685 3582 3418 3598 VDDREF pch l=0.04u w=0.8u
m20686 3587 3419 3599 VDDREF pch l=0.04u w=0.8u
m20687 3586 3421 3601 VDDREF pch l=0.04u w=0.8u
m20688 3622 3422 3602 VDDREF pch l=0.04u w=0.8u
m20689 3589 3423 3603 VDDREF pch l=0.04u w=0.8u
m20690 3588 3425 3605 VDDREF pch l=0.04u w=0.8u
m20691 3623 3426 3606 VDDREF pch l=0.04u w=0.8u
m20692 3782 3708 VDDREF VDDREF pch l=0.04u w=0.8u
m20693 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20694 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m20695 3757 3665 VDDREF VDDREF pch l=0.04u w=0.8u
m20696 3783 3735 VDDREF VDDREF pch l=0.04u w=0.8u
m20697 3768 2508 3180 VDDREF pch l=0.04u w=0.8u
m20698 VDDREF 3835 3764 VDDREF pch l=0.04u w=0.8u
m20699 3765 3953 VDDREF VDDREF pch l=0.04u w=0.8u
m20700 3413 3592 3633 VDDREF pch l=0.04u w=0.8u
m20701 3415 3594 3762 VDDREF pch l=0.04u w=0.8u
m20702 3417 3596 3609 VDDREF pch l=0.04u w=0.8u
m20703 3418 3598 3582 VDDREF pch l=0.04u w=0.8u
m20704 3419 3599 3587 VDDREF pch l=0.04u w=0.8u
m20705 3421 3601 3586 VDDREF pch l=0.04u w=0.8u
m20706 3422 3602 3622 VDDREF pch l=0.04u w=0.8u
m20707 3423 3603 3589 VDDREF pch l=0.04u w=0.8u
m20708 3425 3605 3588 VDDREF pch l=0.04u w=0.8u
m20709 3426 3606 3623 VDDREF pch l=0.04u w=0.8u
m20710 VDDREF 3654 3782 VDDREF pch l=0.04u w=0.8u
m20711 3797 3685 3766 VDDREF pch l=0.04u w=0.8u
m20712 3798 3686 3767 VDDREF pch l=0.04u w=0.8u
m20713 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m20714 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m20715 VDDREF 3849 VDDREF VDDREF pch l=0.26u w=1u
m20716 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20717 3732 3846 VDDREF VDDREF pch l=0.04u w=0.8u
m20718 VDDREF 3713 3757 VDDREF pch l=0.04u w=0.8u
m20719 2508 3180 3768 VDDREF pch l=0.04u w=0.8u
m20720 3799 3680 VDDREF VDDREF pch l=0.04u w=0.8u
m20721 VDDREF 3777 3784 VDDREF pch l=0.04u w=0.8u
m20722 VDDREF 3778 3785 VDDREF pch l=0.04u w=0.8u
m20723 VDDREF 3779 3786 VDDREF pch l=0.04u w=0.8u
m20724 VDDREF 3788 3787 VDDREF pch l=0.04u w=1u
m20725 VDDREF 3789 3790 VDDREF pch l=0.04u w=1u
m20726 VDDREF 3780 3791 VDDREF pch l=0.04u w=0.8u
m20727 VDDREF 3793 3792 VDDREF pch l=0.04u w=1u
m20728 VDDREF 3794 3795 VDDREF pch l=0.04u w=1u
m20729 VDDREF 3781 3796 VDDREF pch l=0.04u w=0.8u
m20730 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20731 31955 4328 3797 VDDREF pch l=0.04u w=0.12u
m20732 31956 4328 3798 VDDREF pch l=0.04u w=0.12u
m20733 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m20734 VDDREF 3867 3732 VDDREF pch l=0.04u w=0.8u
m20735 3800 1200 VDDREF VDDREF pch l=0.04u w=0.8u
m20736 3818 PD VDDREF VDDREF pch l=0.04u w=0.8u
m20737 3819 3694 VDDREF VDDREF pch l=0.04u w=0.8u
m20738 3820 3696 VDDREF VDDREF pch l=0.04u w=0.8u
m20739 3821 3698 VDDREF VDDREF pch l=0.04u w=0.8u
m20740 3822 3699 VDDREF VDDREF pch l=0.04u w=0.8u
m20741 3823 3700 VDDREF VDDREF pch l=0.04u w=0.8u
m20742 3824 3702 VDDREF VDDREF pch l=0.04u w=0.8u
m20743 3825 3703 VDDREF VDDREF pch l=0.04u w=0.8u
m20744 3826 3704 VDDREF VDDREF pch l=0.04u w=0.8u
m20745 3827 3706 VDDREF VDDREF pch l=0.04u w=0.8u
m20746 3828 3707 VDDREF VDDREF pch l=0.04u w=0.8u
m20747 3829 3782 VDDREF VDDREF pch l=0.04u w=0.8u
m20748 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m20749 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m20750 VDDREF 3833 31955 VDDREF pch l=0.04u w=0.12u
m20751 VDDREF 3834 31956 VDDREF pch l=0.04u w=0.12u
m20752 VDDREF 3849 VDDREF VDDREF pch l=0.26u w=1u
m20753 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20754 VDDREF 3801 3802 VDDREF pch l=0.04u w=1u
m20755 VDDREF 3804 3803 VDDREF pch l=0.04u w=1u
m20756 VDDREF 3805 3806 VDDREF pch l=0.04u w=1u
m20757 VDDREF 3808 3807 VDDREF pch l=0.04u w=1u
m20758 VDDREF 3809 3810 VDDREF pch l=0.04u w=1u
m20759 VDDREF 3812 3811 VDDREF pch l=0.04u w=1u
m20760 VDDREF 3813 3814 VDDREF pch l=0.04u w=1u
m20761 VDDREF 3816 3815 VDDREF pch l=0.04u w=1u
m20762 3732 3867 VDDREF VDDREF pch l=0.04u w=0.8u
m20763 3830 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m20764 VDDREF 3906 VDDREF VDDREF pch l=0.26u w=1u
m20765 VDDREF 3907 VDDREF VDDREF pch l=0.26u w=1u
m20766 VDDREF 3910 VDDREF VDDREF pch l=0.26u w=1u
m20767 VDDREF 3911 VDDREF VDDREF pch l=0.26u w=1u
m20768 3817 3768 VDDREF VDDREF pch l=0.04u w=0.8u
m20769 VDDREF 4062 3800 VDDREF pch l=0.04u w=0.8u
m20770 3831 2761 VDDREF VDDREF pch l=0.04u w=0.8u
m20771 3455 3939 VDDREF VDDREF pch l=0.04u w=0.8u
m20772 3457 3940 VDDREF VDDREF pch l=0.04u w=0.8u
m20773 3459 3941 VDDREF VDDREF pch l=0.04u w=0.8u
m20774 3463 3942 VDDREF VDDREF pch l=0.04u w=0.8u
m20775 3467 3943 VDDREF VDDREF pch l=0.04u w=0.8u
m20776 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20777 VDDREF 3727 3829 VDDREF pch l=0.04u w=0.8u
m20778 3833 3797 VDDREF VDDREF pch l=0.04u w=0.8u
m20779 3834 3798 VDDREF VDDREF pch l=0.04u w=0.8u
m20780 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m20781 VDDREF 3846 3732 VDDREF pch l=0.04u w=0.8u
m20782 VDDREF 3666 3817 VDDREF pch l=0.04u w=0.8u
m20783 VDDREF 3025 3831 VDDREF pch l=0.04u w=0.8u
m20784 VDDREF 3854 3455 VDDREF pch l=0.04u w=0.8u
m20785 VDDREF 3855 3457 VDDREF pch l=0.04u w=0.8u
m20786 VDDREF 3856 3459 VDDREF pch l=0.04u w=0.8u
m20787 VDDREF 3857 3463 VDDREF pch l=0.04u w=0.8u
m20788 VDDREF 3858 3467 VDDREF pch l=0.04u w=0.8u
m20789 VDDREF 4251 3832 VDDREF pch l=0.04u w=0.8u
m20790 3836 2780 VDDREF VDDREF pch l=0.04u w=0.8u
m20791 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m20792 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m20793 3837 2781 VDDREF VDDREF pch l=0.04u w=0.8u
m20794 3838 2782 VDDREF VDDREF pch l=0.04u w=0.8u
m20795 3839 2786 VDDREF VDDREF pch l=0.04u w=0.8u
m20796 3840 2787 VDDREF VDDREF pch l=0.04u w=0.8u
m20797 3841 2788 VDDREF VDDREF pch l=0.04u w=0.8u
m20798 3842 2789 VDDREF VDDREF pch l=0.04u w=0.8u
m20799 3843 2790 VDDREF VDDREF pch l=0.04u w=0.8u
m20800 3844 2791 VDDREF VDDREF pch l=0.04u w=0.8u
m20801 3845 2792 VDDREF VDDREF pch l=0.04u w=0.8u
m20802 3829 3727 VDDREF VDDREF pch l=0.04u w=0.8u
m20803 VDDREF 3849 VDDREF VDDREF pch l=0.26u w=1u
m20804 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20805 VDDREF 3921 VDDREF VDDREF pch l=0.26u w=1u
m20806 VDDREF 3924 VDDREF VDDREF pch l=0.26u w=1u
m20807 VDDREF 3925 VDDREF VDDREF pch l=0.26u w=1u
m20808 VDDREF 3928 VDDREF VDDREF pch l=0.26u w=1u
m20809 VDDREF 3929 VDDREF VDDREF pch l=0.26u w=1u
m20810 VDDREF 3932 VDDREF VDDREF pch l=0.26u w=1u
m20811 VDDREF 3933 VDDREF VDDREF pch l=0.26u w=1u
m20812 VDDREF 3936 VDDREF VDDREF pch l=0.26u w=1u
m20813 VDDREF 3906 VDDREF VDDREF pch l=0.26u w=1u
m20814 VDDREF 3907 VDDREF VDDREF pch l=0.26u w=1u
m20815 VDDREF 3910 VDDREF VDDREF pch l=0.26u w=1u
m20816 VDDREF 3911 VDDREF VDDREF pch l=0.26u w=1u
m20817 3847 4251 3757 VDDREF pch l=0.04u w=0.8u
m20818 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20819 3831 3302 VDDREF VDDREF pch l=0.04u w=0.8u
m20820 VDDREF 4062 3835 VDDREF pch l=0.04u w=0.8u
m20821 VDDREF 3047 3836 VDDREF pch l=0.04u w=0.8u
m20822 VDDREF 3049 3837 VDDREF pch l=0.04u w=0.8u
m20823 VDDREF 3051 3838 VDDREF pch l=0.04u w=0.8u
m20824 VDDREF 3053 3839 VDDREF pch l=0.04u w=0.8u
m20825 VDDREF 3054 3840 VDDREF pch l=0.04u w=0.8u
m20826 VDDREF 3056 3841 VDDREF pch l=0.04u w=0.8u
m20827 VDDREF 3057 3842 VDDREF pch l=0.04u w=0.8u
m20828 VDDREF 3058 3843 VDDREF pch l=0.04u w=0.8u
m20829 VDDREF 3060 3844 VDDREF pch l=0.04u w=0.8u
m20830 VDDREF 3061 3845 VDDREF pch l=0.04u w=0.8u
m20831 VDDREF 3782 3829 VDDREF pch l=0.04u w=0.8u
m20832 3848 3848 VDDREF VDDREF pch l=0.04u w=1u
m20833 3850 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20834 3851 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m20835 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m20836 3846 3944 VDDREF VDDREF pch l=0.04u w=0.8u
m20837 31987 3830 3847 VDDREF pch l=0.04u w=0.12u
m20838 3852 3817 VDDREF VDDREF pch l=0.04u w=0.8u
m20839 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m20840 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m20841 3854 3737 VDDREF VDDREF pch l=0.04u w=0.8u
m20842 3836 3321 VDDREF VDDREF pch l=0.04u w=0.8u
m20843 3855 3739 VDDREF VDDREF pch l=0.04u w=0.8u
m20844 3837 3323 VDDREF VDDREF pch l=0.04u w=0.8u
m20845 3856 3741 VDDREF VDDREF pch l=0.04u w=0.8u
m20846 3838 3325 VDDREF VDDREF pch l=0.04u w=0.8u
m20847 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20848 3839 3327 VDDREF VDDREF pch l=0.04u w=0.8u
m20849 3840 3328 VDDREF VDDREF pch l=0.04u w=0.8u
m20850 3857 3745 VDDREF VDDREF pch l=0.04u w=0.8u
m20851 3841 3330 VDDREF VDDREF pch l=0.04u w=0.8u
m20852 3842 3331 VDDREF VDDREF pch l=0.04u w=0.8u
m20853 3843 3332 VDDREF VDDREF pch l=0.04u w=0.8u
m20854 3858 3749 VDDREF VDDREF pch l=0.04u w=0.8u
m20855 3844 3334 VDDREF VDDREF pch l=0.04u w=0.8u
m20856 3845 3335 VDDREF VDDREF pch l=0.04u w=0.8u
m20857 3853 4251 3765 VDDREF pch l=0.04u w=0.8u
m20858 VDDREF 3921 VDDREF VDDREF pch l=0.26u w=1u
m20859 VDDREF 3924 VDDREF VDDREF pch l=0.26u w=1u
m20860 VDDREF 3925 VDDREF VDDREF pch l=0.26u w=1u
m20861 VDDREF 3928 VDDREF VDDREF pch l=0.26u w=1u
m20862 VDDREF 3929 VDDREF VDDREF pch l=0.26u w=1u
m20863 VDDREF 3932 VDDREF VDDREF pch l=0.26u w=1u
m20864 VDDREF 3933 VDDREF VDDREF pch l=0.26u w=1u
m20865 VDDREF 3936 VDDREF VDDREF pch l=0.26u w=1u
m20866 VDDREF 3899 3846 VDDREF pch l=0.04u w=0.8u
m20867 VDDREF 3906 VDDREF VDDREF pch l=0.26u w=1u
m20868 VDDREF 3907 VDDREF VDDREF pch l=0.26u w=1u
m20869 VDDREF 3910 VDDREF VDDREF pch l=0.26u w=1u
m20870 VDDREF 3911 VDDREF VDDREF pch l=0.26u w=1u
m20871 VDDREF 3868 31987 VDDREF pch l=0.04u w=0.12u
m20872 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20873 VDDREF 3714 3852 VDDREF pch l=0.04u w=0.8u
m20874 3861 3831 VDDREF VDDREF pch l=0.04u w=0.8u
m20875 VDDREF 3777 3854 VDDREF pch l=0.04u w=0.8u
m20876 VDDREF 3778 3855 VDDREF pch l=0.04u w=0.8u
m20877 VDDREF 3779 3856 VDDREF pch l=0.04u w=0.8u
m20878 VDDREF 3780 3857 VDDREF pch l=0.04u w=0.8u
m20879 VDDREF 3781 3858 VDDREF pch l=0.04u w=0.8u
m20880 31996 3832 3853 VDDREF pch l=0.04u w=0.12u
m20881 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m20882 3863 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m20883 VDDREF 3860 3859 VDDREF pch l=0.04u w=1u
m20884 3864 4328 3833 VDDREF pch l=0.04u w=0.8u
m20885 3865 4328 3834 VDDREF pch l=0.04u w=0.8u
m20886 3868 3847 VDDREF VDDREF pch l=0.04u w=0.8u
m20887 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m20888 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m20889 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20890 VDDREF 3921 VDDREF VDDREF pch l=0.26u w=1u
m20891 VDDREF 3924 VDDREF VDDREF pch l=0.26u w=1u
m20892 VDDREF 3925 VDDREF VDDREF pch l=0.26u w=1u
m20893 VDDREF 3928 VDDREF VDDREF pch l=0.26u w=1u
m20894 VDDREF 3929 VDDREF VDDREF pch l=0.26u w=1u
m20895 VDDREF 3932 VDDREF VDDREF pch l=0.26u w=1u
m20896 VDDREF 3933 VDDREF VDDREF pch l=0.26u w=1u
m20897 VDDREF 3936 VDDREF VDDREF pch l=0.26u w=1u
m20898 VDDREF 3881 31996 VDDREF pch l=0.04u w=0.12u
m20899 3870 3836 VDDREF VDDREF pch l=0.04u w=0.8u
m20900 3871 3837 VDDREF VDDREF pch l=0.04u w=0.8u
m20901 3872 3838 VDDREF VDDREF pch l=0.04u w=0.8u
m20902 3873 3839 VDDREF VDDREF pch l=0.04u w=0.8u
m20903 3874 3840 VDDREF VDDREF pch l=0.04u w=0.8u
m20904 3875 3841 VDDREF VDDREF pch l=0.04u w=0.8u
m20905 3876 3842 VDDREF VDDREF pch l=0.04u w=0.8u
m20906 3877 3843 VDDREF VDDREF pch l=0.04u w=0.8u
m20907 3878 3844 VDDREF VDDREF pch l=0.04u w=0.8u
m20908 3879 3845 VDDREF VDDREF pch l=0.04u w=0.8u
m20909 3862 3883 3518 VDDREF pch l=0.04u w=0.8u
m20910 32006 3850 3864 VDDREF pch l=0.04u w=0.12u
m20911 32007 3851 3865 VDDREF pch l=0.04u w=0.12u
m20912 VDDREF 3906 VDDREF VDDREF pch l=0.26u w=1u
m20913 VDDREF 3907 VDDREF VDDREF pch l=0.26u w=1u
m20914 VDDREF 3910 VDDREF VDDREF pch l=0.26u w=1u
m20915 VDDREF 3911 VDDREF VDDREF pch l=0.26u w=1u
m20916 3867 FBDIV[9] VDDREF VDDREF pch l=0.04u w=0.8u
m20917 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20918 3880 3768 VDDREF VDDREF pch l=0.04u w=0.8u
m20919 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m20920 3881 3818 VDDREF VDDREF pch l=0.04u w=0.8u
m20921 VDDREF 3968 VDDREF VDDREF pch l=0.26u w=1u
m20922 3882 3861 VDDREF VDDREF pch l=0.04u w=0.8u
m20923 3777 3759 3760 VDDREF pch l=0.04u w=0.8u
m20924 3778 3763 1963 VDDREF pch l=0.04u w=0.8u
m20925 3779 3760 FRAC[12] VDDREF pch l=0.04u w=0.8u
m20926 3780 3553 3409 VDDREF pch l=0.04u w=0.8u
m20927 3781 3554 FRAC[12] VDDREF pch l=0.04u w=0.8u
m20928 3883 3518 3862 VDDREF pch l=0.04u w=0.8u
m20929 3884 4251 3829 VDDREF pch l=0.04u w=0.8u
m20930 VDDREF 3897 32006 VDDREF pch l=0.04u w=0.12u
m20931 VDDREF 3898 32007 VDDREF pch l=0.04u w=0.12u
m20932 VDDREF 4062 3867 VDDREF pch l=0.04u w=0.8u
m20933 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m20934 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m20935 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20936 3885 3830 3868 VDDREF pch l=0.04u w=0.8u
m20937 VDDREF 3921 VDDREF VDDREF pch l=0.26u w=1u
m20938 VDDREF 3924 VDDREF VDDREF pch l=0.26u w=1u
m20939 VDDREF 3925 VDDREF VDDREF pch l=0.26u w=1u
m20940 VDDREF 3928 VDDREF VDDREF pch l=0.26u w=1u
m20941 VDDREF 3929 VDDREF VDDREF pch l=0.26u w=1u
m20942 VDDREF 3932 VDDREF VDDREF pch l=0.26u w=1u
m20943 VDDREF 3933 VDDREF VDDREF pch l=0.26u w=1u
m20944 VDDREF 3936 VDDREF VDDREF pch l=0.26u w=1u
m20945 VDDREF 3853 3881 VDDREF pch l=0.04u w=0.8u
m20946 VDDREF 3569 3882 VDDREF pch l=0.04u w=0.8u
m20947 3759 3760 3777 VDDREF pch l=0.04u w=0.8u
m20948 3763 1963 3778 VDDREF pch l=0.04u w=0.8u
m20949 3760 FRAC[12] 3779 VDDREF pch l=0.04u w=0.8u
m20950 3553 3409 3780 VDDREF pch l=0.04u w=0.8u
m20951 3554 FRAC[12] 3781 VDDREF pch l=0.04u w=0.8u
m20952 VDDREF 3869 3883 VDDREF pch l=0.04u w=0.8u
m20953 3887 3870 VDDREF VDDREF pch l=0.04u w=0.8u
m20954 3888 3871 VDDREF VDDREF pch l=0.04u w=0.8u
m20955 3889 3872 VDDREF VDDREF pch l=0.04u w=0.8u
m20956 3890 3873 VDDREF VDDREF pch l=0.04u w=0.8u
m20957 3891 3874 VDDREF VDDREF pch l=0.04u w=0.8u
m20958 3892 3875 VDDREF VDDREF pch l=0.04u w=0.8u
m20959 3893 3876 VDDREF VDDREF pch l=0.04u w=0.8u
m20960 3894 3877 VDDREF VDDREF pch l=0.04u w=0.8u
m20961 3895 3878 VDDREF VDDREF pch l=0.04u w=0.8u
m20962 3896 3879 VDDREF VDDREF pch l=0.04u w=0.8u
m20963 32024 3863 3884 VDDREF pch l=0.04u w=0.12u
m20964 3897 3864 VDDREF VDDREF pch l=0.04u w=0.8u
m20965 3898 3865 VDDREF VDDREF pch l=0.04u w=0.8u
m20966 VDDREF 3906 VDDREF VDDREF pch l=0.26u w=1u
m20967 VDDREF 3907 VDDREF VDDREF pch l=0.26u w=1u
m20968 VDDREF 3910 VDDREF VDDREF pch l=0.26u w=1u
m20969 VDDREF 3911 VDDREF VDDREF pch l=0.26u w=1u
m20970 VDDREF 3913 VDDREF VDDREF pch l=0.26u w=1u
m20971 32025 4251 3885 VDDREF pch l=0.04u w=0.12u
m20972 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m20973 VDDREF 3968 VDDREF VDDREF pch l=0.26u w=1u
m20974 3886 3666 3768 VDDREF pch l=0.04u w=0.8u
m20975 3882 2667 VDDREF VDDREF pch l=0.04u w=0.8u
m20976 VDDREF 3592 3887 VDDREF pch l=0.04u w=0.8u
m20977 VDDREF 3594 3888 VDDREF pch l=0.04u w=0.8u
m20978 VDDREF 3596 3889 VDDREF pch l=0.04u w=0.8u
m20979 VDDREF 3598 3890 VDDREF pch l=0.04u w=0.8u
m20980 VDDREF 3599 3891 VDDREF pch l=0.04u w=0.8u
m20981 VDDREF 3601 3892 VDDREF pch l=0.04u w=0.8u
m20982 VDDREF 3602 3893 VDDREF pch l=0.04u w=0.8u
m20983 VDDREF 3603 3894 VDDREF pch l=0.04u w=0.8u
m20984 VDDREF 3605 3895 VDDREF pch l=0.04u w=0.8u
m20985 VDDREF 3606 3896 VDDREF pch l=0.04u w=0.8u
m20986 VDDREF 3916 32024 VDDREF pch l=0.04u w=0.12u
m20987 3905 3905 VDDREF VDDREF pch l=0.04u w=1u
m20988 3908 3908 VDDREF VDDREF pch l=0.04u w=1u
m20989 3909 3909 VDDREF VDDREF pch l=0.04u w=1u
m20990 3912 3912 VDDREF VDDREF pch l=0.04u w=1u
m20991 3914 3914 VDDREF VDDREF pch l=0.04u w=1u
m20992 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m20993 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m20994 VDDREF 4062 3899 VDDREF pch l=0.04u w=0.8u
m20995 VDDREF 3920 VDDREF VDDREF pch l=0.26u w=1u
m20996 VDDREF 3921 VDDREF VDDREF pch l=0.26u w=1u
m20997 VDDREF 3924 VDDREF VDDREF pch l=0.26u w=1u
m20998 VDDREF 3925 VDDREF VDDREF pch l=0.26u w=1u
m20999 VDDREF 3928 VDDREF VDDREF pch l=0.26u w=1u
m21000 VDDREF 3929 VDDREF VDDREF pch l=0.26u w=1u
m21001 VDDREF 3932 VDDREF VDDREF pch l=0.26u w=1u
m21002 VDDREF 3933 VDDREF VDDREF pch l=0.26u w=1u
m21003 VDDREF 3936 VDDREF VDDREF pch l=0.26u w=1u
m21004 VDDREF 3590 32025 VDDREF pch l=0.04u w=0.12u
m21005 3666 3768 3886 VDDREF pch l=0.04u w=0.8u
m21006 3915 3832 3881 VDDREF pch l=0.04u w=0.8u
m21007 VDDREF 3759 3900 VDDREF pch l=0.04u w=0.8u
m21008 3887 2678 VDDREF VDDREF pch l=0.04u w=0.8u
m21009 VDDREF 3763 3901 VDDREF pch l=0.04u w=0.8u
m21010 3888 2679 VDDREF VDDREF pch l=0.04u w=0.8u
m21011 VDDREF 3760 3902 VDDREF pch l=0.04u w=0.8u
m21012 3889 2680 VDDREF VDDREF pch l=0.04u w=0.8u
m21013 3890 2683 VDDREF VDDREF pch l=0.04u w=0.8u
m21014 3891 2684 VDDREF VDDREF pch l=0.04u w=0.8u
m21015 VDDREF 3553 3903 VDDREF pch l=0.04u w=0.8u
m21016 3892 2685 VDDREF VDDREF pch l=0.04u w=0.8u
m21017 3893 2686 VDDREF VDDREF pch l=0.04u w=0.8u
m21018 3894 2687 VDDREF VDDREF pch l=0.04u w=0.8u
m21019 VDDREF 3554 3904 VDDREF pch l=0.04u w=0.8u
m21020 3895 2688 VDDREF VDDREF pch l=0.04u w=0.8u
m21021 3896 2689 VDDREF VDDREF pch l=0.04u w=0.8u
m21022 VDDREF 3953 3869 VDDREF pch l=0.04u w=0.8u
m21023 3916 3884 VDDREF VDDREF pch l=0.04u w=0.8u
m21024 3917 3850 3897 VDDREF pch l=0.04u w=0.8u
m21025 3918 3851 3898 VDDREF pch l=0.04u w=0.8u
m21026 3919 3919 VDDREF VDDREF pch l=0.04u w=1u
m21027 3922 3922 VDDREF VDDREF pch l=0.04u w=1u
m21028 3923 3923 VDDREF VDDREF pch l=0.04u w=1u
m21029 3926 3926 VDDREF VDDREF pch l=0.04u w=1u
m21030 3927 3927 VDDREF VDDREF pch l=0.04u w=1u
m21031 3930 3930 VDDREF VDDREF pch l=0.04u w=1u
m21032 3931 3931 VDDREF VDDREF pch l=0.04u w=1u
m21033 3934 3934 VDDREF VDDREF pch l=0.04u w=1u
m21034 3935 3935 VDDREF VDDREF pch l=0.04u w=1u
m21035 VDDREF 3945 VDDREF VDDREF pch l=0.26u w=1u
m21036 3590 3885 VDDREF VDDREF pch l=0.04u w=0.8u
m21037 VDDREF 3968 VDDREF VDDREF pch l=0.26u w=1u
m21038 32042 4251 3915 VDDREF pch l=0.04u w=0.24u
m21039 32043 2445 VDDREF VDDREF pch l=0.04u w=0.8u
m21040 3938 3799 VDDREF VDDREF pch l=0.04u w=0.8u
m21041 32047 4328 3917 VDDREF pch l=0.04u w=0.12u
m21042 32048 4328 3918 VDDREF pch l=0.04u w=0.12u
m21043 VDDREF 3954 VDDREF VDDREF pch l=0.26u w=1u
m21044 VDDREF 3957 VDDREF VDDREF pch l=0.26u w=1u
m21045 3946 3946 VDDREF VDDREF pch l=0.04u w=1u
m21046 VDDREF 4044 32042 VDDREF pch l=0.04u w=0.24u
m21047 3937 3886 32043 VDDREF pch l=0.04u w=0.8u
m21048 VDDREF 3882 3938 VDDREF pch l=0.04u w=0.8u
m21049 3939 3759 VDDREF VDDREF pch l=0.04u w=0.8u
m21050 3737 3819 VDDREF VDDREF pch l=0.04u w=0.8u
m21051 3940 3763 VDDREF VDDREF pch l=0.04u w=0.8u
m21052 3739 3820 VDDREF VDDREF pch l=0.04u w=0.8u
m21053 3941 3760 VDDREF VDDREF pch l=0.04u w=0.8u
m21054 3741 3821 VDDREF VDDREF pch l=0.04u w=0.8u
m21055 3948 3822 VDDREF VDDREF pch l=0.04u w=0.8u
m21056 3949 3823 VDDREF VDDREF pch l=0.04u w=0.8u
m21057 3942 3553 VDDREF VDDREF pch l=0.04u w=0.8u
m21058 3745 3824 VDDREF VDDREF pch l=0.04u w=0.8u
m21059 3950 3825 VDDREF VDDREF pch l=0.04u w=0.8u
m21060 3951 3826 VDDREF VDDREF pch l=0.04u w=0.8u
m21061 3943 3554 VDDREF VDDREF pch l=0.04u w=0.8u
m21062 3749 3827 VDDREF VDDREF pch l=0.04u w=0.8u
m21063 3952 3828 VDDREF VDDREF pch l=0.04u w=0.8u
m21064 3953 3963 VDDREF VDDREF pch l=0.04u w=0.8u
m21065 3947 3863 3916 VDDREF pch l=0.04u w=0.8u
m21066 VDDREF 2131 32047 VDDREF pch l=0.04u w=0.12u
m21067 VDDREF 3961 32048 VDDREF pch l=0.04u w=0.12u
m21068 3955 3955 VDDREF VDDREF pch l=0.04u w=1u
m21069 3956 3956 VDDREF VDDREF pch l=0.04u w=1u
m21070 VDDREF 3968 VDDREF VDDREF pch l=0.26u w=1u
m21071 3944 3962 3619 VDDREF pch l=0.04u w=0.8u
m21072 3959 3590 VDDREF VDDREF pch l=0.04u w=0.8u
m21073 3960 3915 VDDREF VDDREF pch l=0.04u w=0.8u
m21074 VDDREF 3760 3939 VDDREF pch l=0.04u w=0.8u
m21075 VDDREF 3887 3737 VDDREF pch l=0.04u w=0.8u
m21076 VDDREF 1963 3940 VDDREF pch l=0.04u w=0.8u
m21077 VDDREF 3888 3739 VDDREF pch l=0.04u w=0.8u
m21078 VDDREF FRAC[12] 3941 VDDREF pch l=0.04u w=0.8u
m21079 VDDREF 3889 3741 VDDREF pch l=0.04u w=0.8u
m21080 VDDREF 3890 3948 VDDREF pch l=0.04u w=0.8u
m21081 VDDREF 3891 3949 VDDREF pch l=0.04u w=0.8u
m21082 VDDREF 3409 3942 VDDREF pch l=0.04u w=0.8u
m21083 VDDREF 3892 3745 VDDREF pch l=0.04u w=0.8u
m21084 VDDREF 3893 3950 VDDREF pch l=0.04u w=0.8u
m21085 VDDREF 3894 3951 VDDREF pch l=0.04u w=0.8u
m21086 VDDREF FRAC[12] 3943 VDDREF pch l=0.04u w=0.8u
m21087 VDDREF 3895 3749 VDDREF pch l=0.04u w=0.8u
m21088 VDDREF 3896 3952 VDDREF pch l=0.04u w=0.8u
m21089 VDDREF 3963 3953 VDDREF pch l=0.04u w=0.8u
m21090 32069 4251 3947 VDDREF pch l=0.04u w=0.12u
m21091 2131 3917 VDDREF VDDREF pch l=0.04u w=0.8u
m21092 3961 3918 VDDREF VDDREF pch l=0.04u w=0.8u
m21093 3962 3619 3944 VDDREF pch l=0.04u w=0.8u
m21094 VDDREF 3590 3959 VDDREF pch l=0.04u w=0.8u
m21095 VDDREF 3661 32069 VDDREF pch l=0.04u w=0.12u
m21096 VDDREF 3968 VDDREF VDDREF pch l=0.26u w=1u
m21097 VDDREF 3958 3962 VDDREF pch l=0.04u w=0.8u
m21098 3964 3818 VDDREF VDDREF pch l=0.04u w=0.8u
m21099 3661 3947 VDDREF VDDREF pch l=0.04u w=0.8u
m21100 VDDREF 4042 3963 VDDREF pch l=0.04u w=0.8u
m21101 3965 2131 VDDREF VDDREF pch l=0.04u w=0.8u
m21102 3966 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m21103 3967 3967 VDDREF VDDREF pch l=0.04u w=1u
m21104 3969 3959 VDDREF VDDREF pch l=0.04u w=0.8u
m21105 VDDREF 3960 3964 VDDREF pch l=0.04u w=0.8u
m21106 32160 3963 VDDREF VDDREF pch l=0.04u w=0.12u
m21107 3958 3953 VDDREF VDDREF pch l=0.04u w=0.8u
m21108 4042 4251 32160 VDDREF pch l=0.04u w=0.12u
m21109 4040 3661 VDDREF VDDREF pch l=0.04u w=0.8u
m21110 VDDREF 3970 3971 VDDREF pch l=0.04u w=1u
m21111 VDDREF 3973 3972 VDDREF pch l=0.04u w=1u
m21112 VDDREF 3974 3975 VDDREF pch l=0.04u w=1u
m21113 VDDREF 3977 3976 VDDREF pch l=0.04u w=1u
m21114 VDDREF 3978 3979 VDDREF pch l=0.04u w=1u
m21115 VDDREF 3981 3980 VDDREF pch l=0.04u w=1u
m21116 VDDREF 3982 3983 VDDREF pch l=0.04u w=1u
m21117 VDDREF 3985 3984 VDDREF pch l=0.04u w=1u
m21118 VDDREF 3986 3987 VDDREF pch l=0.04u w=1u
m21119 VDDREF 3989 3988 VDDREF pch l=0.04u w=1u
m21120 VDDREF 3990 3991 VDDREF pch l=0.04u w=1u
m21121 VDDREF 3993 3992 VDDREF pch l=0.04u w=1u
m21122 VDDREF 3994 3995 VDDREF pch l=0.04u w=1u
m21123 VDDREF 3997 3996 VDDREF pch l=0.04u w=1u
m21124 VDDREF 3998 3999 VDDREF pch l=0.04u w=1u
m21125 VDDREF 4001 4000 VDDREF pch l=0.04u w=1u
m21126 VDDREF 4002 4003 VDDREF pch l=0.04u w=1u
m21127 VDDREF 4005 4004 VDDREF pch l=0.04u w=1u
m21128 VDDREF 4006 4007 VDDREF pch l=0.04u w=1u
m21129 VDDREF 4009 4008 VDDREF pch l=0.04u w=1u
m21130 4043 4230 VDDREF VDDREF pch l=0.04u w=0.8u
m21131 4041 4328 3961 VDDREF pch l=0.04u w=0.8u
m21132 VDDREF 4010 4011 VDDREF pch l=0.04u w=1u
m21133 VDDREF 4013 4012 VDDREF pch l=0.04u w=1u
m21134 VDDREF 4014 4015 VDDREF pch l=0.04u w=1u
m21135 VDDREF 4017 4016 VDDREF pch l=0.04u w=1u
m21136 VDDREF 4018 4019 VDDREF pch l=0.04u w=1u
m21137 VDDREF 4021 4020 VDDREF pch l=0.04u w=1u
m21138 VDDREF 4022 4023 VDDREF pch l=0.04u w=1u
m21139 VDDREF 4025 4024 VDDREF pch l=0.04u w=1u
m21140 VDDREF 4026 4027 VDDREF pch l=0.04u w=1u
m21141 VDDREF 4029 4028 VDDREF pch l=0.04u w=1u
m21142 VDDREF 4030 4031 VDDREF pch l=0.04u w=1u
m21143 VDDREF 4033 4032 VDDREF pch l=0.04u w=1u
m21144 VDDREF 4034 4035 VDDREF pch l=0.04u w=1u
m21145 VDDREF 4037 4036 VDDREF pch l=0.04u w=1u
m21146 VDDREF 4039 4038 VDDREF pch l=0.04u w=1u
m21147 VDDREF 4048 3958 VDDREF pch l=0.04u w=0.8u
m21148 3567 3524 VDDREF VDDREF pch l=0.04u w=0.8u
m21149 4044 3964 VDDREF VDDREF pch l=0.04u w=0.8u
m21150 4045 4059 4042 VDDREF pch l=0.04u w=0.8u
m21151 VDDREF 3661 4040 VDDREF pch l=0.04u w=0.8u
m21152 32170 3966 4041 VDDREF pch l=0.04u w=0.12u
m21153 4047 4328 VDDREF VDDREF pch l=0.04u w=0.8u
m21154 VDDREF 3969 3567 VDDREF pch l=0.04u w=0.8u
m21155 VDDREF 4068 VDDREF VDDREF pch l=0.26u w=1u
m21156 VDDREF 4071 VDDREF VDDREF pch l=0.26u w=1u
m21157 VDDREF 4072 VDDREF VDDREF pch l=0.26u w=1u
m21158 VDDREF 4075 VDDREF VDDREF pch l=0.26u w=1u
m21159 VDDREF 4076 VDDREF VDDREF pch l=0.26u w=1u
m21160 VDDREF 4079 VDDREF VDDREF pch l=0.26u w=1u
m21161 VDDREF 4080 VDDREF VDDREF pch l=0.26u w=1u
m21162 VDDREF 4083 VDDREF VDDREF pch l=0.26u w=1u
m21163 VDDREF 4084 VDDREF VDDREF pch l=0.26u w=1u
m21164 VDDREF 4087 VDDREF VDDREF pch l=0.26u w=1u
m21165 VDDREF 4088 VDDREF VDDREF pch l=0.26u w=1u
m21166 VDDREF 4091 VDDREF VDDREF pch l=0.26u w=1u
m21167 VDDREF 4092 VDDREF VDDREF pch l=0.26u w=1u
m21168 VDDREF 4095 VDDREF VDDREF pch l=0.26u w=1u
m21169 VDDREF 4096 VDDREF VDDREF pch l=0.26u w=1u
m21170 VDDREF 4099 VDDREF VDDREF pch l=0.26u w=1u
m21171 VDDREF 4100 VDDREF VDDREF pch l=0.26u w=1u
m21172 VDDREF 4103 VDDREF VDDREF pch l=0.26u w=1u
m21173 VDDREF 4104 VDDREF VDDREF pch l=0.26u w=1u
m21174 VDDREF 4107 VDDREF VDDREF pch l=0.26u w=1u
m21175 VDDREF 4108 VDDREF VDDREF pch l=0.26u w=1u
m21176 VDDREF 4111 VDDREF VDDREF pch l=0.26u w=1u
m21177 VDDREF 4112 VDDREF VDDREF pch l=0.26u w=1u
m21178 VDDREF 4115 VDDREF VDDREF pch l=0.26u w=1u
m21179 VDDREF 4116 VDDREF VDDREF pch l=0.26u w=1u
m21180 VDDREF 4119 VDDREF VDDREF pch l=0.26u w=1u
m21181 VDDREF 4120 VDDREF VDDREF pch l=0.26u w=1u
m21182 VDDREF 4123 VDDREF VDDREF pch l=0.26u w=1u
m21183 VDDREF 4124 VDDREF VDDREF pch l=0.26u w=1u
m21184 VDDREF 4127 VDDREF VDDREF pch l=0.26u w=1u
m21185 VDDREF 4128 VDDREF VDDREF pch l=0.26u w=1u
m21186 VDDREF 4131 VDDREF VDDREF pch l=0.26u w=1u
m21187 VDDREF 4132 VDDREF VDDREF pch l=0.26u w=1u
m21188 VDDREF 4135 VDDREF VDDREF pch l=0.26u w=1u
m21189 VDDREF 4051 32170 VDDREF pch l=0.04u w=0.12u
m21190 VDDREF 4328 4046 VDDREF pch l=0.04u w=0.8u
m21191 VDDREF 4139 VDDREF VDDREF pch l=0.26u w=1u
m21192 VDDREF 4053 4048 VDDREF pch l=0.04u w=0.8u
m21193 4049 3964 VDDREF VDDREF pch l=0.04u w=0.8u
m21194 VDDREF 4057 4045 VDDREF pch l=0.04u w=0.8u
m21195 4050 4040 VDDREF VDDREF pch l=0.04u w=0.8u
m21196 4051 4041 VDDREF VDDREF pch l=0.04u w=0.8u
m21197 CLKSSCG 4047 VDDREF VDDREF pch l=0.04u w=0.8u
m21198 4054 3524 VDDREF VDDREF pch l=0.04u w=0.8u
m21199 VDDREF 4068 VDDREF VDDREF pch l=0.26u w=1u
m21200 VDDREF 4071 VDDREF VDDREF pch l=0.26u w=1u
m21201 VDDREF 4072 VDDREF VDDREF pch l=0.26u w=1u
m21202 VDDREF 4075 VDDREF VDDREF pch l=0.26u w=1u
m21203 VDDREF 4076 VDDREF VDDREF pch l=0.26u w=1u
m21204 VDDREF 4079 VDDREF VDDREF pch l=0.26u w=1u
m21205 VDDREF 4080 VDDREF VDDREF pch l=0.26u w=1u
m21206 VDDREF 4083 VDDREF VDDREF pch l=0.26u w=1u
m21207 VDDREF 4084 VDDREF VDDREF pch l=0.26u w=1u
m21208 VDDREF 4087 VDDREF VDDREF pch l=0.26u w=1u
m21209 VDDREF 4088 VDDREF VDDREF pch l=0.26u w=1u
m21210 VDDREF 4091 VDDREF VDDREF pch l=0.26u w=1u
m21211 VDDREF 4092 VDDREF VDDREF pch l=0.26u w=1u
m21212 VDDREF 4095 VDDREF VDDREF pch l=0.26u w=1u
m21213 VDDREF 4096 VDDREF VDDREF pch l=0.26u w=1u
m21214 VDDREF 4099 VDDREF VDDREF pch l=0.26u w=1u
m21215 VDDREF 4100 VDDREF VDDREF pch l=0.26u w=1u
m21216 VDDREF 4103 VDDREF VDDREF pch l=0.26u w=1u
m21217 VDDREF 4104 VDDREF VDDREF pch l=0.26u w=1u
m21218 VDDREF 4107 VDDREF VDDREF pch l=0.26u w=1u
m21219 VDDREF 4108 VDDREF VDDREF pch l=0.26u w=1u
m21220 VDDREF 4111 VDDREF VDDREF pch l=0.26u w=1u
m21221 VDDREF 4112 VDDREF VDDREF pch l=0.26u w=1u
m21222 VDDREF 4115 VDDREF VDDREF pch l=0.26u w=1u
m21223 VDDREF 4116 VDDREF VDDREF pch l=0.26u w=1u
m21224 VDDREF 4119 VDDREF VDDREF pch l=0.26u w=1u
m21225 VDDREF 4120 VDDREF VDDREF pch l=0.26u w=1u
m21226 VDDREF 4123 VDDREF VDDREF pch l=0.26u w=1u
m21227 VDDREF 4124 VDDREF VDDREF pch l=0.26u w=1u
m21228 VDDREF 4127 VDDREF VDDREF pch l=0.26u w=1u
m21229 VDDREF 4128 VDDREF VDDREF pch l=0.26u w=1u
m21230 VDDREF 4131 VDDREF VDDREF pch l=0.26u w=1u
m21231 VDDREF 4132 VDDREF VDDREF pch l=0.26u w=1u
m21232 VDDREF 4135 VDDREF VDDREF pch l=0.26u w=1u
m21233 VDDREF 3964 4049 VDDREF pch l=0.04u w=0.8u
m21234 32188 4045 VDDREF VDDREF pch l=0.04u w=0.12u
m21235 VDDREF 3450 4050 VDDREF pch l=0.04u w=0.8u
m21236 VDDREF 4139 VDDREF VDDREF pch l=0.26u w=1u
m21237 4055 4328 3965 VDDREF pch l=0.04u w=0.8u
m21238 VDDREF 4047 CLKSSCG VDDREF pch l=0.04u w=0.8u
m21239 VDDREF 3484 4053 VDDREF pch l=0.04u w=0.8u
m21240 VDDREF 3959 4054 VDDREF pch l=0.04u w=0.8u
m21241 4049 3964 VDDREF VDDREF pch l=0.04u w=0.8u
m21242 4057 4059 32188 VDDREF pch l=0.04u w=0.12u
m21243 4050 2969 VDDREF VDDREF pch l=0.04u w=0.8u
m21244 4056 3966 4051 VDDREF pch l=0.04u w=0.8u
m21245 32193 4046 4055 VDDREF pch l=0.04u w=0.12u
m21246 CLKSSCG 4047 VDDREF VDDREF pch l=0.04u w=0.8u
m21247 4053 4351 VDDREF VDDREF pch l=0.04u w=0.8u
m21248 4054 3959 VDDREF VDDREF pch l=0.04u w=0.8u
m21249 VDDREF 4068 VDDREF VDDREF pch l=0.26u w=1u
m21250 VDDREF 4071 VDDREF VDDREF pch l=0.26u w=1u
m21251 VDDREF 4072 VDDREF VDDREF pch l=0.26u w=1u
m21252 VDDREF 4075 VDDREF VDDREF pch l=0.26u w=1u
m21253 VDDREF 4076 VDDREF VDDREF pch l=0.26u w=1u
m21254 VDDREF 4079 VDDREF VDDREF pch l=0.26u w=1u
m21255 VDDREF 4080 VDDREF VDDREF pch l=0.26u w=1u
m21256 VDDREF 4083 VDDREF VDDREF pch l=0.26u w=1u
m21257 VDDREF 4084 VDDREF VDDREF pch l=0.26u w=1u
m21258 VDDREF 4087 VDDREF VDDREF pch l=0.26u w=1u
m21259 VDDREF 4088 VDDREF VDDREF pch l=0.26u w=1u
m21260 VDDREF 4091 VDDREF VDDREF pch l=0.26u w=1u
m21261 VDDREF 4092 VDDREF VDDREF pch l=0.26u w=1u
m21262 VDDREF 4095 VDDREF VDDREF pch l=0.26u w=1u
m21263 VDDREF 4096 VDDREF VDDREF pch l=0.26u w=1u
m21264 VDDREF 4099 VDDREF VDDREF pch l=0.26u w=1u
m21265 VDDREF 4100 VDDREF VDDREF pch l=0.26u w=1u
m21266 VDDREF 4103 VDDREF VDDREF pch l=0.26u w=1u
m21267 VDDREF 4104 VDDREF VDDREF pch l=0.26u w=1u
m21268 VDDREF 4107 VDDREF VDDREF pch l=0.26u w=1u
m21269 VDDREF 4108 VDDREF VDDREF pch l=0.26u w=1u
m21270 VDDREF 4111 VDDREF VDDREF pch l=0.26u w=1u
m21271 VDDREF 4112 VDDREF VDDREF pch l=0.26u w=1u
m21272 VDDREF 4115 VDDREF VDDREF pch l=0.26u w=1u
m21273 VDDREF 4116 VDDREF VDDREF pch l=0.26u w=1u
m21274 VDDREF 4119 VDDREF VDDREF pch l=0.26u w=1u
m21275 VDDREF 4120 VDDREF VDDREF pch l=0.26u w=1u
m21276 VDDREF 4123 VDDREF VDDREF pch l=0.26u w=1u
m21277 VDDREF 4124 VDDREF VDDREF pch l=0.26u w=1u
m21278 VDDREF 4127 VDDREF VDDREF pch l=0.26u w=1u
m21279 VDDREF 4128 VDDREF VDDREF pch l=0.26u w=1u
m21280 VDDREF 4131 VDDREF VDDREF pch l=0.26u w=1u
m21281 VDDREF 4132 VDDREF VDDREF pch l=0.26u w=1u
m21282 VDDREF 4135 VDDREF VDDREF pch l=0.26u w=1u
m21283 VDDREF 3964 4049 VDDREF pch l=0.04u w=0.8u
m21284 4058 4251 4057 VDDREF pch l=0.04u w=0.8u
m21285 VDDREF 4139 VDDREF VDDREF pch l=0.26u w=1u
m21286 32201 4328 4056 VDDREF pch l=0.04u w=0.12u
m21287 VDDREF 4061 32193 VDDREF pch l=0.04u w=0.12u
m21288 VDDREF 4047 CLKSSCG VDDREF pch l=0.04u w=0.8u
m21289 VDDREF 4064 4053 VDDREF pch l=0.04u w=0.8u
m21290 VDDREF 3524 4054 VDDREF pch l=0.04u w=0.8u
m21291 4060 4050 VDDREF VDDREF pch l=0.04u w=0.8u
m21292 VDDREF 4063 32201 VDDREF pch l=0.04u w=0.12u
m21293 4061 4043 VDDREF VDDREF pch l=0.04u w=0.8u
m21294 VDDREF 4068 VDDREF VDDREF pch l=0.26u w=1u
m21295 VDDREF 4071 VDDREF VDDREF pch l=0.26u w=1u
m21296 VDDREF 4072 VDDREF VDDREF pch l=0.26u w=1u
m21297 VDDREF 4075 VDDREF VDDREF pch l=0.26u w=1u
m21298 VDDREF 4076 VDDREF VDDREF pch l=0.26u w=1u
m21299 VDDREF 4079 VDDREF VDDREF pch l=0.26u w=1u
m21300 VDDREF 4080 VDDREF VDDREF pch l=0.26u w=1u
m21301 VDDREF 4083 VDDREF VDDREF pch l=0.26u w=1u
m21302 VDDREF 4084 VDDREF VDDREF pch l=0.26u w=1u
m21303 VDDREF 4087 VDDREF VDDREF pch l=0.26u w=1u
m21304 VDDREF 4088 VDDREF VDDREF pch l=0.26u w=1u
m21305 VDDREF 4091 VDDREF VDDREF pch l=0.26u w=1u
m21306 VDDREF 4092 VDDREF VDDREF pch l=0.26u w=1u
m21307 VDDREF 4095 VDDREF VDDREF pch l=0.26u w=1u
m21308 VDDREF 4096 VDDREF VDDREF pch l=0.26u w=1u
m21309 VDDREF 4099 VDDREF VDDREF pch l=0.26u w=1u
m21310 VDDREF 4100 VDDREF VDDREF pch l=0.26u w=1u
m21311 VDDREF 4103 VDDREF VDDREF pch l=0.26u w=1u
m21312 VDDREF 4104 VDDREF VDDREF pch l=0.26u w=1u
m21313 VDDREF 4107 VDDREF VDDREF pch l=0.26u w=1u
m21314 VDDREF 4108 VDDREF VDDREF pch l=0.26u w=1u
m21315 VDDREF 4111 VDDREF VDDREF pch l=0.26u w=1u
m21316 VDDREF 4112 VDDREF VDDREF pch l=0.26u w=1u
m21317 VDDREF 4115 VDDREF VDDREF pch l=0.26u w=1u
m21318 VDDREF 4116 VDDREF VDDREF pch l=0.26u w=1u
m21319 VDDREF 4119 VDDREF VDDREF pch l=0.26u w=1u
m21320 VDDREF 4120 VDDREF VDDREF pch l=0.26u w=1u
m21321 VDDREF 4123 VDDREF VDDREF pch l=0.26u w=1u
m21322 VDDREF 4124 VDDREF VDDREF pch l=0.26u w=1u
m21323 VDDREF 4127 VDDREF VDDREF pch l=0.26u w=1u
m21324 VDDREF 4128 VDDREF VDDREF pch l=0.26u w=1u
m21325 VDDREF 4131 VDDREF VDDREF pch l=0.26u w=1u
m21326 VDDREF 4132 VDDREF VDDREF pch l=0.26u w=1u
m21327 VDDREF 4135 VDDREF VDDREF pch l=0.26u w=1u
m21328 4062 4049 VDDREF VDDREF pch l=0.04u w=0.8u
m21329 VDDREF 4139 VDDREF VDDREF pch l=0.26u w=1u
m21330 VDDREF 4251 4059 VDDREF pch l=0.04u w=0.8u
m21331 4063 4056 VDDREF VDDREF pch l=0.04u w=0.8u
m21332 VDDREF 4055 4061 VDDREF pch l=0.04u w=0.8u
m21333 4064 4136 VDDREF VDDREF pch l=0.04u w=0.8u
m21334 3117 4054 VDDREF VDDREF pch l=0.04u w=0.8u
m21335 VDDREF 4049 4062 VDDREF pch l=0.04u w=0.8u
m21336 4065 4060 VDDREF VDDREF pch l=0.04u w=0.8u
m21337 VDDREF 4068 VDDREF VDDREF pch l=0.26u w=1u
m21338 VDDREF 4071 VDDREF VDDREF pch l=0.26u w=1u
m21339 VDDREF 4072 VDDREF VDDREF pch l=0.26u w=1u
m21340 VDDREF 4075 VDDREF VDDREF pch l=0.26u w=1u
m21341 VDDREF 4076 VDDREF VDDREF pch l=0.26u w=1u
m21342 VDDREF 4079 VDDREF VDDREF pch l=0.26u w=1u
m21343 VDDREF 4080 VDDREF VDDREF pch l=0.26u w=1u
m21344 VDDREF 4083 VDDREF VDDREF pch l=0.26u w=1u
m21345 VDDREF 4084 VDDREF VDDREF pch l=0.26u w=1u
m21346 VDDREF 4087 VDDREF VDDREF pch l=0.26u w=1u
m21347 VDDREF 4088 VDDREF VDDREF pch l=0.26u w=1u
m21348 VDDREF 4091 VDDREF VDDREF pch l=0.26u w=1u
m21349 VDDREF 4092 VDDREF VDDREF pch l=0.26u w=1u
m21350 VDDREF 4095 VDDREF VDDREF pch l=0.26u w=1u
m21351 VDDREF 4096 VDDREF VDDREF pch l=0.26u w=1u
m21352 VDDREF 4099 VDDREF VDDREF pch l=0.26u w=1u
m21353 VDDREF 4100 VDDREF VDDREF pch l=0.26u w=1u
m21354 VDDREF 4103 VDDREF VDDREF pch l=0.26u w=1u
m21355 VDDREF 4104 VDDREF VDDREF pch l=0.26u w=1u
m21356 VDDREF 4107 VDDREF VDDREF pch l=0.26u w=1u
m21357 VDDREF 4108 VDDREF VDDREF pch l=0.26u w=1u
m21358 VDDREF 4111 VDDREF VDDREF pch l=0.26u w=1u
m21359 VDDREF 4112 VDDREF VDDREF pch l=0.26u w=1u
m21360 VDDREF 4115 VDDREF VDDREF pch l=0.26u w=1u
m21361 VDDREF 4116 VDDREF VDDREF pch l=0.26u w=1u
m21362 VDDREF 4119 VDDREF VDDREF pch l=0.26u w=1u
m21363 VDDREF 4120 VDDREF VDDREF pch l=0.26u w=1u
m21364 VDDREF 4123 VDDREF VDDREF pch l=0.26u w=1u
m21365 VDDREF 4124 VDDREF VDDREF pch l=0.26u w=1u
m21366 VDDREF 4127 VDDREF VDDREF pch l=0.26u w=1u
m21367 VDDREF 4128 VDDREF VDDREF pch l=0.26u w=1u
m21368 VDDREF 4131 VDDREF VDDREF pch l=0.26u w=1u
m21369 VDDREF 4132 VDDREF VDDREF pch l=0.26u w=1u
m21370 VDDREF 4135 VDDREF VDDREF pch l=0.26u w=1u
m21371 VDDREF 4136 4064 VDDREF pch l=0.04u w=0.8u
m21372 VDDREF 4139 VDDREF VDDREF pch l=0.26u w=1u
m21373 4062 4049 VDDREF VDDREF pch l=0.04u w=0.8u
m21374 4058 4218 VDDREF VDDREF pch l=0.04u w=0.8u
m21375 VDDREF 3484 4065 VDDREF pch l=0.04u w=0.8u
m21376 4067 4063 VDDREF VDDREF pch l=0.04u w=0.8u
m21377 4066 4046 4061 VDDREF pch l=0.04u w=0.8u
m21378 4069 4069 VDDREF VDDREF pch l=0.04u w=1u
m21379 4070 4070 VDDREF VDDREF pch l=0.04u w=1u
m21380 4073 4073 VDDREF VDDREF pch l=0.04u w=1u
m21381 4074 4074 VDDREF VDDREF pch l=0.04u w=1u
m21382 4077 4077 VDDREF VDDREF pch l=0.04u w=1u
m21383 4078 4078 VDDREF VDDREF pch l=0.04u w=1u
m21384 4081 4081 VDDREF VDDREF pch l=0.04u w=1u
m21385 4082 4082 VDDREF VDDREF pch l=0.04u w=1u
m21386 4085 4085 VDDREF VDDREF pch l=0.04u w=1u
m21387 4086 4086 VDDREF VDDREF pch l=0.04u w=1u
m21388 4089 4089 VDDREF VDDREF pch l=0.04u w=1u
m21389 4090 4090 VDDREF VDDREF pch l=0.04u w=1u
m21390 4093 4093 VDDREF VDDREF pch l=0.04u w=1u
m21391 4094 4094 VDDREF VDDREF pch l=0.04u w=1u
m21392 4097 4097 VDDREF VDDREF pch l=0.04u w=1u
m21393 4098 4098 VDDREF VDDREF pch l=0.04u w=1u
m21394 4101 4101 VDDREF VDDREF pch l=0.04u w=1u
m21395 4102 4102 VDDREF VDDREF pch l=0.04u w=1u
m21396 4105 4105 VDDREF VDDREF pch l=0.04u w=1u
m21397 4106 4106 VDDREF VDDREF pch l=0.04u w=1u
m21398 4109 4109 VDDREF VDDREF pch l=0.04u w=1u
m21399 4110 4110 VDDREF VDDREF pch l=0.04u w=1u
m21400 4113 4113 VDDREF VDDREF pch l=0.04u w=1u
m21401 4114 4114 VDDREF VDDREF pch l=0.04u w=1u
m21402 4117 4117 VDDREF VDDREF pch l=0.04u w=1u
m21403 4118 4118 VDDREF VDDREF pch l=0.04u w=1u
m21404 4121 4121 VDDREF VDDREF pch l=0.04u w=1u
m21405 4122 4122 VDDREF VDDREF pch l=0.04u w=1u
m21406 4125 4125 VDDREF VDDREF pch l=0.04u w=1u
m21407 4126 4126 VDDREF VDDREF pch l=0.04u w=1u
m21408 4129 4129 VDDREF VDDREF pch l=0.04u w=1u
m21409 4130 4130 VDDREF VDDREF pch l=0.04u w=1u
m21410 4133 4133 VDDREF VDDREF pch l=0.04u w=1u
m21411 4134 4134 VDDREF VDDREF pch l=0.04u w=1u
m21412 4137 4363 VDDREF VDDREF pch l=0.04u w=0.8u
m21413 4138 4138 VDDREF VDDREF pch l=0.04u w=1u
m21414 VDDREF 4049 4062 VDDREF pch l=0.04u w=0.8u
m21415 VDDREF 4224 4058 VDDREF pch l=0.04u w=0.8u
m21416 4065 3953 VDDREF VDDREF pch l=0.04u w=0.8u
m21417 32234 4328 4066 VDDREF pch l=0.04u w=0.24u
m21418 VDDREF 4216 4136 VDDREF pch l=0.04u w=0.8u
m21419 VDDREF 4054 4137 VDDREF pch l=0.04u w=0.8u
m21420 4062 4049 VDDREF VDDREF pch l=0.04u w=0.8u
m21421 4058 4224 VDDREF VDDREF pch l=0.04u w=0.8u
m21422 VDDREF 4226 32234 VDDREF pch l=0.04u w=0.24u
m21423 4212 4230 VDDREF VDDREF pch l=0.04u w=0.8u
m21424 VDDREF 4140 4141 VDDREF pch l=0.04u w=1u
m21425 VDDREF 4143 4142 VDDREF pch l=0.04u w=1u
m21426 VDDREF 4144 4145 VDDREF pch l=0.04u w=1u
m21427 VDDREF 4147 4146 VDDREF pch l=0.04u w=1u
m21428 VDDREF 4148 4149 VDDREF pch l=0.04u w=1u
m21429 VDDREF 4151 4150 VDDREF pch l=0.04u w=1u
m21430 VDDREF 4152 4153 VDDREF pch l=0.04u w=1u
m21431 VDDREF 4155 4154 VDDREF pch l=0.04u w=1u
m21432 VDDREF 4156 4157 VDDREF pch l=0.04u w=1u
m21433 VDDREF 4159 4158 VDDREF pch l=0.04u w=1u
m21434 VDDREF 4160 4161 VDDREF pch l=0.04u w=1u
m21435 VDDREF 4163 4162 VDDREF pch l=0.04u w=1u
m21436 VDDREF 4164 4165 VDDREF pch l=0.04u w=1u
m21437 VDDREF 4167 4166 VDDREF pch l=0.04u w=1u
m21438 VDDREF 4168 4169 VDDREF pch l=0.04u w=1u
m21439 VDDREF 4171 4170 VDDREF pch l=0.04u w=1u
m21440 VDDREF 4172 4173 VDDREF pch l=0.04u w=1u
m21441 VDDREF 4175 4174 VDDREF pch l=0.04u w=1u
m21442 VDDREF 4176 4177 VDDREF pch l=0.04u w=1u
m21443 VDDREF 4179 4178 VDDREF pch l=0.04u w=1u
m21444 VDDREF 4180 4181 VDDREF pch l=0.04u w=1u
m21445 VDDREF 4183 4182 VDDREF pch l=0.04u w=1u
m21446 VDDREF 4184 4185 VDDREF pch l=0.04u w=1u
m21447 VDDREF 4187 4186 VDDREF pch l=0.04u w=1u
m21448 VDDREF 4188 4189 VDDREF pch l=0.04u w=1u
m21449 VDDREF 4191 4190 VDDREF pch l=0.04u w=1u
m21450 VDDREF 4192 4193 VDDREF pch l=0.04u w=1u
m21451 VDDREF 4195 4194 VDDREF pch l=0.04u w=1u
m21452 VDDREF 4196 4197 VDDREF pch l=0.04u w=1u
m21453 VDDREF 4199 4198 VDDREF pch l=0.04u w=1u
m21454 VDDREF 4200 4201 VDDREF pch l=0.04u w=1u
m21455 VDDREF 4203 4202 VDDREF pch l=0.04u w=1u
m21456 VDDREF 4204 4205 VDDREF pch l=0.04u w=1u
m21457 VDDREF 4207 4206 VDDREF pch l=0.04u w=1u
m21458 VDDREF 4208 4209 VDDREF pch l=0.04u w=1u
m21459 32242 4136 VDDREF VDDREF pch l=0.04u w=0.12u
m21460 VDDREF 4049 4062 VDDREF pch l=0.04u w=0.8u
m21461 VDDREF 4211 4210 VDDREF pch l=0.04u w=1u
m21462 VDDREF 4218 4058 VDDREF pch l=0.04u w=0.8u
m21463 4213 4065 VDDREF VDDREF pch l=0.04u w=0.8u
m21464 4214 4066 VDDREF VDDREF pch l=0.04u w=0.8u
m21465 4216 4251 32242 VDDREF pch l=0.04u w=0.12u
m21466 4217 4617 VDDREF VDDREF pch l=0.04u w=0.8u
m21467 4219 4221 4213 VDDREF pch l=0.04u w=0.8u
m21468 VDDREF 4328 4215 VDDREF pch l=0.04u w=0.8u
m21469 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21470 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21471 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21472 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21473 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21474 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21475 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21476 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21477 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21478 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21479 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21480 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21481 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21482 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21483 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21484 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21485 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21486 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21487 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21488 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21489 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21490 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21491 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21492 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21493 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21494 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21495 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21496 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21497 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21498 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21499 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21500 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21501 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21502 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21503 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21504 4220 4234 4216 VDDREF pch l=0.04u w=0.8u
m21505 VDDREF 4241 VDDREF VDDREF pch l=0.26u w=1u
m21506 4062 4049 VDDREF VDDREF pch l=0.04u w=0.8u
m21507 4218 4238 VDDREF VDDREF pch l=0.04u w=0.8u
m21508 4221 4213 4219 VDDREF pch l=0.04u w=0.8u
m21509 69 4043 VDDREF VDDREF pch l=0.04u w=0.8u
m21510 4222 4617 4137 VDDREF pch l=0.04u w=0.8u
m21511 VDDREF 4049 4062 VDDREF pch l=0.04u w=0.8u
m21512 VDDREF 4232 4218 VDDREF pch l=0.04u w=0.8u
m21513 VDDREF 4214 69 VDDREF pch l=0.04u w=0.8u
m21514 4223 4328 4067 VDDREF pch l=0.04u w=0.8u
m21515 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21516 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21517 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21518 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21519 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21520 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21521 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21522 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21523 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21524 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21525 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21526 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21527 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21528 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21529 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21530 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21531 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21532 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21533 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21534 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21535 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21536 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21537 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21538 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21539 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21540 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21541 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21542 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21543 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21544 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21545 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21546 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21547 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21548 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21549 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21550 VDDREF 4241 VDDREF VDDREF pch l=0.26u w=1u
m21551 VDDREF 4227 4220 VDDREF pch l=0.04u w=0.8u
m21552 32265 4217 4222 VDDREF pch l=0.04u w=0.12u
m21553 4062 4049 VDDREF VDDREF pch l=0.04u w=0.8u
m21554 32267 4215 4223 VDDREF pch l=0.04u w=0.12u
m21555 32274 4220 VDDREF VDDREF pch l=0.04u w=0.12u
m21556 VDDREF 4228 32265 VDDREF pch l=0.04u w=0.12u
m21557 VDDREF 4049 4062 VDDREF pch l=0.04u w=0.8u
m21558 4224 911 VDDREF VDDREF pch l=0.04u w=0.8u
m21559 4225 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m21560 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21561 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21562 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21563 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21564 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21565 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21566 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21567 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21568 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21569 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21570 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21571 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21572 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21573 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21574 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21575 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21576 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21577 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21578 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21579 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21580 4226 69 VDDREF VDDREF pch l=0.04u w=0.8u
m21581 VDDREF 4229 32267 VDDREF pch l=0.04u w=0.12u
m21582 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21583 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21584 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21585 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21586 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21587 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21588 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21589 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21590 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21591 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21592 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21593 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21594 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21595 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21596 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21597 VDDREF 4241 VDDREF VDDREF pch l=0.26u w=1u
m21598 4227 4234 32274 VDDREF pch l=0.04u w=0.12u
m21599 4228 4222 VDDREF VDDREF pch l=0.04u w=0.8u
m21600 4062 4049 VDDREF VDDREF pch l=0.04u w=0.8u
m21601 VDDREF 4062 4224 VDDREF pch l=0.04u w=0.8u
m21602 4229 4212 VDDREF VDDREF pch l=0.04u w=0.8u
m21603 4231 4251 4227 VDDREF pch l=0.04u w=0.8u
m21604 VDDREF 4049 4062 VDDREF pch l=0.04u w=0.8u
m21605 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21606 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21607 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21608 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21609 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21610 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21611 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21612 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21613 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21614 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21615 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21616 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21617 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21618 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21619 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21620 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21621 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21622 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21623 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21624 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21625 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21626 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21627 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21628 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21629 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21630 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21631 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21632 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21633 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21634 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21635 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21636 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21637 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21638 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21639 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21640 VDDREF 4223 4229 VDDREF pch l=0.04u w=0.8u
m21641 4233 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m21642 VDDREF 2616 4230 VDDREF pch l=0.04u w=0.8u
m21643 VDDREF 4241 VDDREF VDDREF pch l=0.26u w=1u
m21644 4235 4217 4228 VDDREF pch l=0.04u w=0.8u
m21645 VDDREF 4062 4232 VDDREF pch l=0.04u w=0.8u
m21646 VDDREF 2501 4233 VDDREF pch l=0.04u w=0.8u
m21647 VDDREF 4251 4234 VDDREF pch l=0.04u w=0.8u
m21648 32297 4617 4235 VDDREF pch l=0.04u w=0.12u
m21649 4236 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m21650 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21651 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21652 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21653 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21654 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21655 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21656 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21657 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21658 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21659 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21660 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21661 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21662 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21663 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21664 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21665 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21666 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21667 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21668 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21669 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21670 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21671 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21672 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21673 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21674 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21675 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21676 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21677 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21678 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21679 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21680 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21681 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21682 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21683 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21684 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21685 4237 4215 4229 VDDREF pch l=0.04u w=0.8u
m21686 VDDREF 4241 VDDREF VDDREF pch l=0.26u w=1u
m21687 VDDREF 4242 32297 VDDREF pch l=0.04u w=0.12u
m21688 32310 4328 4237 VDDREF pch l=0.04u w=0.24u
m21689 4239 4225 VDDREF VDDREF pch l=0.04u w=0.8u
m21690 4240 4240 VDDREF VDDREF pch l=0.04u w=1u
m21691 4231 4250 VDDREF VDDREF pch l=0.04u w=0.8u
m21692 4242 4235 VDDREF VDDREF pch l=0.04u w=0.8u
m21693 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21694 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21695 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21696 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21697 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21698 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21699 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21700 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21701 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21702 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21703 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21704 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21705 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21706 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21707 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21708 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21709 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21710 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21711 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21712 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21713 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21714 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21715 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21716 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21717 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21718 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21719 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21720 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21721 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21722 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21723 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21724 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21725 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21726 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21727 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21728 4243 4251 4062 VDDREF pch l=0.04u w=0.8u
m21729 VDDREF 4324 32310 VDDREF pch l=0.04u w=0.24u
m21730 4238 4245 3963 VDDREF pch l=0.04u w=0.8u
m21731 VDDREF 4219 4239 VDDREF pch l=0.04u w=0.8u
m21732 VDDREF 4325 4231 VDDREF pch l=0.04u w=0.8u
m21733 32350 4236 4243 VDDREF pch l=0.04u w=0.12u
m21734 4244 4237 VDDREF VDDREF pch l=0.04u w=0.8u
m21735 4245 3963 4238 VDDREF pch l=0.04u w=0.8u
m21736 4231 4325 VDDREF VDDREF pch l=0.04u w=0.8u
m21737 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21738 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21739 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21740 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21741 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21742 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21743 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21744 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21745 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21746 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21747 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21748 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21749 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21750 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21751 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21752 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21753 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21754 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21755 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21756 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21757 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21758 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21759 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21760 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21761 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21762 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21763 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21764 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21765 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21766 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21767 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21768 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21769 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21770 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21771 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21772 4246 4242 VDDREF VDDREF pch l=0.04u w=0.8u
m21773 VDDREF 4249 32350 VDDREF pch l=0.04u w=0.12u
m21774 VDDREF PD 4245 VDDREF pch l=0.04u w=0.8u
m21775 4247 4239 VDDREF VDDREF pch l=0.04u w=0.8u
m21776 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21777 VDDREF 4250 4231 VDDREF pch l=0.04u w=0.8u
m21778 VDDREF 4359 4246 VDDREF pch l=0.04u w=0.8u
m21779 4249 4243 VDDREF VDDREF pch l=0.04u w=0.8u
m21780 70 4212 VDDREF VDDREF pch l=0.04u w=0.8u
m21781 VDDREF 4233 4247 VDDREF pch l=0.04u w=0.8u
m21782 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21783 VDDREF 4252 VDDREF VDDREF pch l=0.26u w=1u
m21784 VDDREF 4255 VDDREF VDDREF pch l=0.26u w=1u
m21785 VDDREF 4256 VDDREF VDDREF pch l=0.26u w=1u
m21786 VDDREF 4259 VDDREF VDDREF pch l=0.26u w=1u
m21787 VDDREF 4260 VDDREF VDDREF pch l=0.26u w=1u
m21788 VDDREF 4263 VDDREF VDDREF pch l=0.26u w=1u
m21789 VDDREF 4264 VDDREF VDDREF pch l=0.26u w=1u
m21790 VDDREF 4267 VDDREF VDDREF pch l=0.26u w=1u
m21791 VDDREF 4268 VDDREF VDDREF pch l=0.26u w=1u
m21792 VDDREF 4271 VDDREF VDDREF pch l=0.26u w=1u
m21793 VDDREF 4272 VDDREF VDDREF pch l=0.26u w=1u
m21794 VDDREF 4275 VDDREF VDDREF pch l=0.26u w=1u
m21795 VDDREF 4276 VDDREF VDDREF pch l=0.26u w=1u
m21796 VDDREF 4279 VDDREF VDDREF pch l=0.26u w=1u
m21797 VDDREF 4280 VDDREF VDDREF pch l=0.26u w=1u
m21798 VDDREF 4283 VDDREF VDDREF pch l=0.26u w=1u
m21799 VDDREF 4284 VDDREF VDDREF pch l=0.26u w=1u
m21800 VDDREF 4287 VDDREF VDDREF pch l=0.26u w=1u
m21801 VDDREF 4288 VDDREF VDDREF pch l=0.26u w=1u
m21802 VDDREF 4291 VDDREF VDDREF pch l=0.26u w=1u
m21803 VDDREF 4292 VDDREF VDDREF pch l=0.26u w=1u
m21804 VDDREF 4295 VDDREF VDDREF pch l=0.26u w=1u
m21805 VDDREF 4296 VDDREF VDDREF pch l=0.26u w=1u
m21806 VDDREF 4299 VDDREF VDDREF pch l=0.26u w=1u
m21807 VDDREF 4300 VDDREF VDDREF pch l=0.26u w=1u
m21808 VDDREF 4303 VDDREF VDDREF pch l=0.26u w=1u
m21809 VDDREF 4304 VDDREF VDDREF pch l=0.26u w=1u
m21810 VDDREF 4307 VDDREF VDDREF pch l=0.26u w=1u
m21811 VDDREF 4308 VDDREF VDDREF pch l=0.26u w=1u
m21812 VDDREF 4311 VDDREF VDDREF pch l=0.26u w=1u
m21813 VDDREF 4312 VDDREF VDDREF pch l=0.26u w=1u
m21814 VDDREF 4315 VDDREF VDDREF pch l=0.26u w=1u
m21815 VDDREF 4316 VDDREF VDDREF pch l=0.26u w=1u
m21816 VDDREF 4319 VDDREF VDDREF pch l=0.26u w=1u
m21817 VDDREF 4320 VDDREF VDDREF pch l=0.26u w=1u
m21818 VDDREF 4244 70 VDDREF pch l=0.04u w=0.8u
m21819 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21820 4247 4233 VDDREF VDDREF pch l=0.04u w=0.8u
m21821 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21822 4253 4253 VDDREF VDDREF pch l=0.04u w=1u
m21823 4254 4254 VDDREF VDDREF pch l=0.04u w=1u
m21824 4257 4257 VDDREF VDDREF pch l=0.04u w=1u
m21825 4258 4258 VDDREF VDDREF pch l=0.04u w=1u
m21826 4261 4261 VDDREF VDDREF pch l=0.04u w=1u
m21827 4262 4262 VDDREF VDDREF pch l=0.04u w=1u
m21828 4265 4265 VDDREF VDDREF pch l=0.04u w=1u
m21829 4266 4266 VDDREF VDDREF pch l=0.04u w=1u
m21830 4269 4269 VDDREF VDDREF pch l=0.04u w=1u
m21831 4270 4270 VDDREF VDDREF pch l=0.04u w=1u
m21832 4273 4273 VDDREF VDDREF pch l=0.04u w=1u
m21833 4274 4274 VDDREF VDDREF pch l=0.04u w=1u
m21834 4277 4277 VDDREF VDDREF pch l=0.04u w=1u
m21835 4278 4278 VDDREF VDDREF pch l=0.04u w=1u
m21836 4281 4281 VDDREF VDDREF pch l=0.04u w=1u
m21837 4282 4282 VDDREF VDDREF pch l=0.04u w=1u
m21838 4285 4285 VDDREF VDDREF pch l=0.04u w=1u
m21839 4286 4286 VDDREF VDDREF pch l=0.04u w=1u
m21840 4289 4289 VDDREF VDDREF pch l=0.04u w=1u
m21841 4290 4290 VDDREF VDDREF pch l=0.04u w=1u
m21842 4293 4293 VDDREF VDDREF pch l=0.04u w=1u
m21843 4294 4294 VDDREF VDDREF pch l=0.04u w=1u
m21844 4297 4297 VDDREF VDDREF pch l=0.04u w=1u
m21845 4298 4298 VDDREF VDDREF pch l=0.04u w=1u
m21846 4301 4301 VDDREF VDDREF pch l=0.04u w=1u
m21847 4302 4302 VDDREF VDDREF pch l=0.04u w=1u
m21848 4305 4305 VDDREF VDDREF pch l=0.04u w=1u
m21849 4306 4306 VDDREF VDDREF pch l=0.04u w=1u
m21850 4309 4309 VDDREF VDDREF pch l=0.04u w=1u
m21851 4310 4310 VDDREF VDDREF pch l=0.04u w=1u
m21852 4313 4313 VDDREF VDDREF pch l=0.04u w=1u
m21853 4314 4314 VDDREF VDDREF pch l=0.04u w=1u
m21854 4317 4317 VDDREF VDDREF pch l=0.04u w=1u
m21855 4318 4318 VDDREF VDDREF pch l=0.04u w=1u
m21856 4321 4321 VDDREF VDDREF pch l=0.04u w=1u
m21857 4250 4337 VDDREF VDDREF pch l=0.04u w=0.8u
m21858 4322 4617 VDDREF VDDREF pch l=0.04u w=0.8u
m21859 4323 4249 VDDREF VDDREF pch l=0.04u w=0.8u
m21860 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21861 VDDREF 4239 4247 VDDREF pch l=0.04u w=0.8u
m21862 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21863 VDDREF 4331 4250 VDDREF pch l=0.04u w=0.8u
m21864 VDDREF 4249 4323 VDDREF pch l=0.04u w=0.8u
m21865 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21866 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21867 4324 70 VDDREF VDDREF pch l=0.04u w=0.8u
m21868 4326 4617 4246 VDDREF pch l=0.04u w=0.8u
m21869 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21870 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21871 4327 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m21872 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21873 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21874 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21875 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21876 4325 2952 VDDREF VDDREF pch l=0.04u w=0.8u
m21877 32499 4322 4326 VDDREF pch l=0.04u w=0.12u
m21878 4329 4062 VDDREF VDDREF pch l=0.04u w=0.8u
m21879 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21880 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21881 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21882 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21883 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21884 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21885 VDDREF 4062 4325 VDDREF pch l=0.04u w=0.8u
m21886 VDDREF 4332 32499 VDDREF pch l=0.04u w=0.12u
m21887 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21888 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21889 4330 4251 4247 VDDREF pch l=0.04u w=0.8u
m21890 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21891 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21892 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21893 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21894 4332 4326 VDDREF VDDREF pch l=0.04u w=0.8u
m21895 4333 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m21896 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21897 32773 4327 4330 VDDREF pch l=0.04u w=0.12u
m21898 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21899 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21900 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21901 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21902 VDDREF 4062 4331 VDDREF pch l=0.04u w=0.8u
m21903 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21904 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21905 VDDREF 4336 32773 VDDREF pch l=0.04u w=0.12u
m21906 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21907 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21908 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21909 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21910 4334 4322 4332 VDDREF pch l=0.04u w=0.8u
m21911 4335 4251 4329 VDDREF pch l=0.04u w=0.8u
m21912 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21913 4336 4330 VDDREF VDDREF pch l=0.04u w=0.8u
m21914 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21915 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21916 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21917 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21918 33141 4617 4334 VDDREF pch l=0.04u w=0.12u
m21919 33142 4333 4335 VDDREF pch l=0.04u w=0.12u
m21920 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21921 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21922 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21923 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21924 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21925 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21926 VDDREF 4340 33141 VDDREF pch l=0.04u w=0.12u
m21927 4337 4341 4136 VDDREF pch l=0.04u w=0.8u
m21928 VDDREF 4342 33142 VDDREF pch l=0.04u w=0.12u
m21929 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21930 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21931 4339 4327 4336 VDDREF pch l=0.04u w=0.8u
m21932 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21933 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21934 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21935 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21936 4340 4334 VDDREF VDDREF pch l=0.04u w=0.8u
m21937 4341 4136 4337 VDDREF pch l=0.04u w=0.8u
m21938 4342 4335 VDDREF VDDREF pch l=0.04u w=0.8u
m21939 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21940 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21941 33698 4251 4339 VDDREF pch l=0.04u w=0.12u
m21942 VDDREF 4338 4341 VDDREF pch l=0.04u w=0.8u
m21943 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21944 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21945 VDDREF 4221 33698 VDDREF pch l=0.04u w=0.12u
m21946 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21947 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21948 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21949 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21950 4343 4617 VDDREF VDDREF pch l=0.04u w=0.8u
m21951 4344 4333 4342 VDDREF pch l=0.04u w=0.8u
m21952 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21953 4248 4346 VDDREF VDDREF pch l=0.04u w=0.8u
m21954 4221 4339 VDDREF VDDREF pch l=0.04u w=0.8u
m21955 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21956 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21957 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21958 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21959 VDDREF 3953 4338 VDDREF pch l=0.04u w=0.8u
m21960 34068 4251 4344 VDDREF pch l=0.04u w=0.12u
m21961 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21962 VDDREF 4346 4248 VDDREF pch l=0.04u w=0.8u
m21963 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21964 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21965 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21966 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21967 4338 3484 VDDREF VDDREF pch l=0.04u w=0.8u
m21968 4345 4617 4340 VDDREF pch l=0.04u w=0.8u
m21969 VDDREF 4348 34068 VDDREF pch l=0.04u w=0.12u
m21970 4251 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21971 4347 4221 VDDREF VDDREF pch l=0.04u w=0.8u
m21972 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21973 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21974 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21975 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21976 VDDREF 4351 4338 VDDREF pch l=0.04u w=0.8u
m21977 34437 4343 4345 VDDREF pch l=0.04u w=0.12u
m21978 4348 4344 VDDREF VDDREF pch l=0.04u w=0.8u
m21979 VDDREF 4362 4251 VDDREF pch l=0.04u w=0.8u
m21980 VDDREF 4368 4346 VDDREF pch l=0.04u w=0.4u
m21981 VDDREF 4221 4347 VDDREF pch l=0.04u w=0.8u
m21982 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21983 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21984 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21985 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21986 VDDREF 4350 34437 VDDREF pch l=0.04u w=0.12u
m21987 4346 4368 VDDREF VDDREF pch l=0.04u w=0.4u
m21988 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21989 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21990 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21991 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m21992 4350 4345 VDDREF VDDREF pch l=0.04u w=0.8u
m21993 4351 4357 VDDREF VDDREF pch l=0.04u w=0.8u
m21994 4352 4251 VDDREF VDDREF pch l=0.04u w=0.8u
m21995 4353 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m21996 VDDREF 4368 4346 VDDREF pch l=0.04u w=0.4u
m21997 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21998 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m21999 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m22000 4328 4248 VDDREF VDDREF pch l=0.04u w=0.8u
m22001 VDDREF 4357 4351 VDDREF pch l=0.04u w=0.8u
m22002 VDDREF 4362 4353 VDDREF pch l=0.04u w=0.8u
m22003 4346 4368 VDDREF VDDREF pch l=0.04u w=0.4u
m22004 VDDREF 4354 4355 VDDREF pch l=0.04u w=1u
m22005 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m22006 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m22007 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m22008 VDDREF 4248 4328 VDDREF pch l=0.04u w=0.8u
m22009 4356 4343 4350 VDDREF pch l=0.04u w=0.8u
m22010 4353 4362 VDDREF VDDREF pch l=0.04u w=0.8u
m22011 4358 4251 4348 VDDREF pch l=0.04u w=0.8u
m22012 VDDREF 4368 4346 VDDREF pch l=0.04u w=0.4u
m22013 34664 4617 4356 VDDREF pch l=0.04u w=0.12u
m22014 4357 2969 VDDREF VDDREF pch l=0.04u w=0.8u
m22015 VDDREF 4362 4353 VDDREF pch l=0.04u w=0.8u
m22016 34665 4352 4358 VDDREF pch l=0.04u w=0.12u
m22017 4346 4368 VDDREF VDDREF pch l=0.04u w=0.4u
m22018 VDDREF 4369 VDDREF VDDREF pch l=0.26u w=1u
m22019 VDDREF 4359 34664 VDDREF pch l=0.04u w=0.12u
m22020 VDDREF 4360 4357 VDDREF pch l=0.04u w=0.8u
m22021 VDDREF 4361 34665 VDDREF pch l=0.04u w=0.12u
m22022 VDDREF 4368 4346 VDDREF pch l=0.04u w=0.4u
m22023 4359 4356 VDDREF VDDREF pch l=0.04u w=0.8u
m22024 4361 4358 VDDREF VDDREF pch l=0.04u w=0.8u
m22025 4346 4368 VDDREF VDDREF pch l=0.04u w=0.4u
m22026 4362 4366 VDDREF VDDREF pch l=0.04u w=0.8u
m22027 VDDREF 4369 VDDREF VDDREF pch l=0.26u w=1u
m22028 VDDREF 4365 4360 VDDREF pch l=0.04u w=0.8u
m22029 VDDREF 4367 4346 VDDREF pch l=0.04u w=0.4u
m22030 VDDREF 4366 4362 VDDREF pch l=0.04u w=0.8u
m22031 4363 4359 VDDREF VDDREF pch l=0.04u w=0.8u
m22032 4362 4366 VDDREF VDDREF pch l=0.04u w=0.8u
m22033 VDDREF 4369 VDDREF VDDREF pch l=0.26u w=1u
m22034 4364 4352 4361 VDDREF pch l=0.04u w=0.8u
m22035 VDDREF 4366 4362 VDDREF pch l=0.04u w=0.8u
m22036 VDDREF 3450 4365 VDDREF pch l=0.04u w=0.8u
m22037 34744 4251 4364 VDDREF pch l=0.04u w=0.12u
m22038 VDDREF 4369 VDDREF VDDREF pch l=0.26u w=1u
m22039 4366 4363 VDDREF VDDREF pch l=0.04u w=0.8u
m22040 4362 4366 VDDREF VDDREF pch l=0.04u w=0.8u
m22041 4365 4040 VDDREF VDDREF pch l=0.04u w=0.8u
m22042 VDDREF 4368 34744 VDDREF pch l=0.04u w=0.12u
m22043 VDDREF 4363 4366 VDDREF pch l=0.04u w=0.8u
m22044 VDDREF 4366 4362 VDDREF pch l=0.04u w=0.8u
m22045 VDDREF 4347 4365 VDDREF pch l=0.04u w=0.8u
m22046 4368 4364 VDDREF VDDREF pch l=0.04u w=0.8u
m22047 VDDREF DSMPD 4367 VDDREF pch l=0.04u w=0.8u
m22048 VDDREF 4369 VDDREF VDDREF pch l=0.26u w=1u
m22049 4370 4370 VDDREF VDDREF pch l=0.04u w=1u
m22050 VDDREF 4372 4371 VDDREF pch l=0.04u w=1u
m22051 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22052 VDDPOST 4374 4375 VDDPOST pch l=0.04u w=1u
m22053 VDDPOST 4377 4376 VDDPOST pch l=0.04u w=1u
m22054 VDDREF 4378 4379 VDDREF pch l=0.04u w=1u
m22055 VDDREF 4381 4380 VDDREF pch l=0.04u w=1u
m22056 VDDREF 4382 4383 VDDREF pch l=0.04u w=1u
m22057 VDDREF 4385 4384 VDDREF pch l=0.04u w=1u
m22058 VDDREF 4386 4387 VDDREF pch l=0.04u w=1u
m22059 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22060 4388 2427 VDDREF VDDREF pch l=0.04u w=0.8u
m22061 4390 4390 VDDREF VDDREF pch l=0.04u w=1u
m22062 VDDREF 2427 4388 VDDREF pch l=0.04u w=0.8u
m22063 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22064 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22065 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22066 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22067 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22068 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22069 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22070 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22071 34956 FBDIV[10] VDDREF VDDREF pch l=0.04u w=0.8u
m22072 4392 2426 VDDREF VDDREF pch l=0.04u w=0.8u
m22073 4391 FBDIV[11] 34956 VDDREF pch l=0.04u w=0.8u
m22074 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22075 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22076 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22077 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22078 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22079 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22080 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22081 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22082 VDDREF 2426 4392 VDDREF pch l=0.04u w=0.8u
m22083 34980 2952 VDDREF VDDREF pch l=0.04u w=0.8u
m22084 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22085 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22086 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22087 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22088 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22089 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22090 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22091 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22092 4394 4323 VDDREF VDDREF pch l=0.04u w=0.8u
m22093 4393 FBDIV[9] 34980 VDDREF pch l=0.04u w=0.8u
m22094 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22095 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22096 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22097 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22098 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22099 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22100 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22101 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22102 4395 4394 VDDREF VDDREF pch l=0.04u w=0.8u
m22103 4396 4393 VDDREF VDDREF pch l=0.04u w=0.8u
m22104 VDDREF 4394 4395 VDDREF pch l=0.04u w=0.8u
m22105 VDDREF 4391 4396 VDDREF pch l=0.04u w=0.8u
m22106 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22107 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22108 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22109 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22110 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22111 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22112 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22113 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22114 4395 4394 VDDREF VDDREF pch l=0.04u w=0.8u
m22115 VDDREF 4394 4395 VDDREF pch l=0.04u w=0.8u
m22116 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22117 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22118 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22119 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22120 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22121 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22122 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22123 4397 2427 VDDREF VDDREF pch l=0.04u w=0.8u
m22124 VDDREF 4399 VDDREF VDDREF pch l=0.26u w=1u
m22125 4398 4398 VDDREF VDDREF pch l=0.04u w=1u
m22126 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22127 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22128 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22129 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22130 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22131 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22132 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22133 35565 3293 VDDREF VDDREF pch l=0.04u w=0.8u
m22134 4401 DSMPD VDDREF VDDREF pch l=0.04u w=0.8u
m22135 4400 3783 35565 VDDREF pch l=0.04u w=0.8u
m22136 VDDREF 4396 4401 VDDREF pch l=0.04u w=0.8u
m22137 VDDREF 4403 4402 VDDREF pch l=0.04u w=1u
m22138 VDDPOST 4404 VDDPOST VDDPOST pch l=0.26u w=1u
m22139 VDDPOST 4407 VDDPOST VDDPOST pch l=0.26u w=1u
m22140 VDDREF 4408 VDDREF VDDREF pch l=0.26u w=1u
m22141 VDDREF 4411 VDDREF VDDREF pch l=0.26u w=1u
m22142 VDDREF 4412 VDDREF VDDREF pch l=0.26u w=1u
m22143 VDDREF 4415 VDDREF VDDREF pch l=0.26u w=1u
m22144 VDDREF 4416 VDDREF VDDREF pch l=0.26u w=1u
m22145 4401 4397 VDDREF VDDREF pch l=0.04u w=0.8u
m22146 4405 4405 VDDPOST VDDPOST pch l=0.04u w=1u
m22147 4406 4406 VDDPOST VDDPOST pch l=0.04u w=1u
m22148 4409 4409 VDDREF VDDREF pch l=0.04u w=1u
m22149 4410 4410 VDDREF VDDREF pch l=0.04u w=1u
m22150 4413 4413 VDDREF VDDREF pch l=0.04u w=1u
m22151 4414 4414 VDDREF VDDREF pch l=0.04u w=1u
m22152 4417 4417 VDDREF VDDREF pch l=0.04u w=1u
m22153 4418 4400 VDDREF VDDREF pch l=0.04u w=0.8u
m22154 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22155 4423 DSMPD VDDREF VDDREF pch l=0.04u w=0.8u
m22156 VDDPOST 4419 4420 VDDPOST pch l=0.04u w=1u
m22157 VDDPOST 4422 4421 VDDPOST pch l=0.04u w=1u
m22158 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22159 35828 3480 VDDREF VDDREF pch l=0.04u w=0.8u
m22160 VDDREF 4396 4423 VDDREF pch l=0.04u w=0.8u
m22161 4424 3937 35828 VDDREF pch l=0.04u w=0.8u
m22162 4423 2426 VDDREF VDDREF pch l=0.04u w=0.8u
m22163 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22164 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22165 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22166 4425 4424 VDDREF VDDREF pch l=0.04u w=0.8u
m22167 4426 4423 VDDREF VDDREF pch l=0.04u w=0.8u
m22168 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22169 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22170 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22171 4427 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22172 4428 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22173 4429 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22174 4430 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22175 4431 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22176 4432 4467 VDDREF VDDREF pch l=0.04u w=0.8u
m22177 4433 4468 VDDREF VDDREF pch l=0.04u w=0.8u
m22178 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22179 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22180 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22181 VDDREF 2509 4427 VDDREF pch l=0.04u w=0.8u
m22182 VDDREF 2747 4428 VDDREF pch l=0.04u w=0.8u
m22183 VDDREF 3019 4429 VDDREF pch l=0.04u w=0.8u
m22184 VDDREF 4418 4430 VDDREF pch l=0.04u w=0.8u
m22185 VDDREF 3783 4431 VDDREF pch l=0.04u w=0.8u
m22186 VDDREF 4467 4432 VDDREF pch l=0.04u w=0.8u
m22187 VDDREF 4468 4433 VDDREF pch l=0.04u w=0.8u
m22188 4432 4467 VDDREF VDDREF pch l=0.04u w=0.8u
m22189 4433 4468 VDDREF VDDREF pch l=0.04u w=0.8u
m22190 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22191 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22192 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22193 VDDREF 4467 4432 VDDREF pch l=0.04u w=0.8u
m22194 VDDREF 4468 4433 VDDREF pch l=0.04u w=0.8u
m22195 4434 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22196 4435 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22197 4436 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22198 4437 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22199 4438 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22200 4432 4467 VDDREF VDDREF pch l=0.04u w=0.8u
m22201 4433 4468 VDDREF VDDREF pch l=0.04u w=0.8u
m22202 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22203 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22204 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22205 VDDREF 4467 4432 VDDREF pch l=0.04u w=0.8u
m22206 VDDREF 4468 4433 VDDREF pch l=0.04u w=0.8u
m22207 4439 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22208 4440 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22209 4441 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22210 4442 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22211 4443 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22212 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22213 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22214 VDDREF DACPD 4439 VDDREF pch l=0.04u w=0.8u
m22215 VDDREF DACPD 4440 VDDREF pch l=0.04u w=0.8u
m22216 VDDREF DACPD 4441 VDDREF pch l=0.04u w=0.8u
m22217 VDDREF DACPD 4442 VDDREF pch l=0.04u w=0.8u
m22218 VDDREF DACPD 4443 VDDREF pch l=0.04u w=0.8u
m22219 VDDREF 4446 VDDREF VDDREF pch l=0.26u w=1u
m22220 4432 4467 VDDREF VDDREF pch l=0.04u w=0.8u
m22221 4433 4468 VDDREF VDDREF pch l=0.04u w=0.8u
m22222 4445 4445 VDDREF VDDREF pch l=0.04u w=1u
m22223 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22224 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22225 VDDREF 4467 4432 VDDREF pch l=0.04u w=0.8u
m22226 VDDREF 4468 4433 VDDREF pch l=0.04u w=0.8u
m22227 4447 4434 VDDREF VDDREF pch l=0.04u w=0.8u
m22228 4448 4435 VDDREF VDDREF pch l=0.04u w=0.8u
m22229 4449 4436 VDDREF VDDREF pch l=0.04u w=0.8u
m22230 4450 4437 VDDREF VDDREF pch l=0.04u w=0.8u
m22231 4451 4438 VDDREF VDDREF pch l=0.04u w=0.8u
m22232 4432 4467 VDDREF VDDREF pch l=0.04u w=0.8u
m22233 4433 4468 VDDREF VDDREF pch l=0.04u w=0.8u
m22234 VDDREF 4427 4447 VDDREF pch l=0.04u w=0.8u
m22235 VDDREF 4428 4448 VDDREF pch l=0.04u w=0.8u
m22236 VDDREF 4429 4449 VDDREF pch l=0.04u w=0.8u
m22237 VDDREF 4430 4450 VDDREF pch l=0.04u w=0.8u
m22238 VDDREF 4431 4451 VDDREF pch l=0.04u w=0.8u
m22239 VDDREF 4453 4452 VDDREF pch l=0.04u w=1u
m22240 VDDPOST 4454 VDDPOST VDDPOST pch l=0.26u w=1u
m22241 VDDPOST 4457 VDDPOST VDDPOST pch l=0.26u w=1u
m22242 VDDREF 4467 4432 VDDREF pch l=0.04u w=0.8u
m22243 VDDREF 4468 4433 VDDREF pch l=0.04u w=0.8u
m22244 4455 4455 VDDPOST VDDPOST pch l=0.04u w=1u
m22245 4456 4456 VDDPOST VDDPOST pch l=0.04u w=1u
m22246 4432 4467 VDDREF VDDREF pch l=0.04u w=0.8u
m22247 4433 4468 VDDREF VDDREF pch l=0.04u w=0.8u
m22248 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22249 4458 4447 VDDREF VDDREF pch l=0.04u w=0.8u
m22250 4459 4448 VDDREF VDDREF pch l=0.04u w=0.8u
m22251 4460 4449 VDDREF VDDREF pch l=0.04u w=0.8u
m22252 4461 4450 VDDREF VDDREF pch l=0.04u w=0.8u
m22253 4462 4451 VDDREF VDDREF pch l=0.04u w=0.8u
m22254 VDDREF 4467 4432 VDDREF pch l=0.04u w=0.8u
m22255 VDDREF 4468 4433 VDDREF pch l=0.04u w=0.8u
m22256 VDDREF 4439 4458 VDDREF pch l=0.04u w=0.8u
m22257 VDDREF 4440 4459 VDDREF pch l=0.04u w=0.8u
m22258 VDDREF 4441 4460 VDDREF pch l=0.04u w=0.8u
m22259 VDDREF 4442 4461 VDDREF pch l=0.04u w=0.8u
m22260 VDDREF 4443 4462 VDDREF pch l=0.04u w=0.8u
m22261 VDDPOST 4463 4464 VDDPOST pch l=0.04u w=1u
m22262 VDDPOST 4466 4465 VDDPOST pch l=0.04u w=1u
m22263 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22264 4467 4480 VDDREF VDDREF pch l=0.04u w=0.8u
m22265 4468 4481 VDDREF VDDREF pch l=0.04u w=0.8u
m22266 4469 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22267 4470 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22268 4471 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22269 4472 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22270 4473 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22271 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22272 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22273 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22274 VDDREF 4480 4467 VDDREF pch l=0.04u w=0.8u
m22275 VDDREF 4481 4468 VDDREF pch l=0.04u w=0.8u
m22276 4467 4480 VDDREF VDDREF pch l=0.04u w=0.8u
m22277 4468 4481 VDDREF VDDREF pch l=0.04u w=0.8u
m22278 4475 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22279 4476 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22280 4477 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22281 4478 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22282 4479 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22283 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22284 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22285 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22286 VDDREF 4480 4467 VDDREF pch l=0.04u w=0.8u
m22287 VDDREF 4481 4468 VDDREF pch l=0.04u w=0.8u
m22288 VDDREF 4388 4475 VDDREF pch l=0.04u w=0.8u
m22289 VDDREF 4388 4476 VDDREF pch l=0.04u w=0.8u
m22290 VDDREF 4388 4477 VDDREF pch l=0.04u w=0.8u
m22291 VDDREF 4388 4478 VDDREF pch l=0.04u w=0.8u
m22292 VDDREF 4388 4479 VDDREF pch l=0.04u w=0.8u
m22293 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22294 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22295 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22296 4480 4502 VDDREF VDDREF pch l=0.04u w=0.8u
m22297 4481 4503 VDDREF VDDREF pch l=0.04u w=0.8u
m22298 4482 4469 VDDREF VDDREF pch l=0.04u w=0.8u
m22299 4483 4470 VDDREF VDDREF pch l=0.04u w=0.8u
m22300 4484 4471 VDDREF VDDREF pch l=0.04u w=0.8u
m22301 4485 4472 VDDREF VDDREF pch l=0.04u w=0.8u
m22302 4486 4473 VDDREF VDDREF pch l=0.04u w=0.8u
m22303 VDDREF 2427 4480 VDDREF pch l=0.04u w=0.8u
m22304 VDDREF 4401 4481 VDDREF pch l=0.04u w=0.8u
m22305 VDDREF 4458 4482 VDDREF pch l=0.04u w=0.8u
m22306 VDDREF 4459 4483 VDDREF pch l=0.04u w=0.8u
m22307 VDDREF 4460 4484 VDDREF pch l=0.04u w=0.8u
m22308 VDDREF 4461 4485 VDDREF pch l=0.04u w=0.8u
m22309 VDDREF 4462 4486 VDDREF pch l=0.04u w=0.8u
m22310 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22311 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22312 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22313 4480 2427 VDDREF VDDREF pch l=0.04u w=0.8u
m22314 4481 4401 VDDREF VDDREF pch l=0.04u w=0.8u
m22315 VDDREF 4502 4480 VDDREF pch l=0.04u w=0.8u
m22316 VDDREF 4503 4481 VDDREF pch l=0.04u w=0.8u
m22317 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22318 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22319 4487 4482 VDDREF VDDREF pch l=0.04u w=0.8u
m22320 4488 4483 VDDREF VDDREF pch l=0.04u w=0.8u
m22321 4489 4484 VDDREF VDDREF pch l=0.04u w=0.8u
m22322 4490 4485 VDDREF VDDREF pch l=0.04u w=0.8u
m22323 4491 4486 VDDREF VDDREF pch l=0.04u w=0.8u
m22324 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22325 VDDREF 4475 4487 VDDREF pch l=0.04u w=0.8u
m22326 VDDREF 4476 4488 VDDREF pch l=0.04u w=0.8u
m22327 VDDREF 4477 4489 VDDREF pch l=0.04u w=0.8u
m22328 VDDREF 4478 4490 VDDREF pch l=0.04u w=0.8u
m22329 VDDREF 4479 4491 VDDREF pch l=0.04u w=0.8u
m22330 4493 2427 VDDREF VDDREF pch l=0.04u w=0.8u
m22331 4494 4401 VDDREF VDDREF pch l=0.04u w=0.8u
m22332 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22333 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22334 VDDREF 4496 VDDREF VDDREF pch l=0.26u w=1u
m22335 4495 4495 VDDREF VDDREF pch l=0.04u w=1u
m22336 4497 4487 VDDREF VDDREF pch l=0.04u w=0.8u
m22337 4498 4488 VDDREF VDDREF pch l=0.04u w=0.8u
m22338 4499 4489 VDDREF VDDREF pch l=0.04u w=0.8u
m22339 4500 4490 VDDREF VDDREF pch l=0.04u w=0.8u
m22340 4501 4491 VDDREF VDDREF pch l=0.04u w=0.8u
m22341 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22342 4502 4480 VDDREF VDDREF pch l=0.04u w=0.8u
m22343 4503 4481 VDDREF VDDREF pch l=0.04u w=0.8u
m22344 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22345 VDDREF 4493 4502 VDDREF pch l=0.04u w=0.8u
m22346 VDDREF 4494 4503 VDDREF pch l=0.04u w=0.8u
m22347 VDDREF 4505 4504 VDDREF pch l=0.04u w=1u
m22348 4506 4522 VDDREF VDDREF pch l=0.04u w=0.8u
m22349 4507 4523 VDDREF VDDREF pch l=0.04u w=0.8u
m22350 4508 4524 VDDREF VDDREF pch l=0.04u w=0.8u
m22351 4509 4525 VDDREF VDDREF pch l=0.04u w=0.8u
m22352 4510 4526 VDDREF VDDREF pch l=0.04u w=0.8u
m22353 VDDPOST 4511 VDDPOST VDDPOST pch l=0.26u w=1u
m22354 VDDPOST 4514 VDDPOST VDDPOST pch l=0.26u w=1u
m22355 4502 4493 VDDREF VDDREF pch l=0.04u w=0.8u
m22356 4503 4494 VDDREF VDDREF pch l=0.04u w=0.8u
m22357 VDDREF 4522 4506 VDDREF pch l=0.04u w=0.8u
m22358 VDDREF 4523 4507 VDDREF pch l=0.04u w=0.8u
m22359 VDDREF 4524 4508 VDDREF pch l=0.04u w=0.8u
m22360 VDDREF 4525 4509 VDDREF pch l=0.04u w=0.8u
m22361 VDDREF 4526 4510 VDDREF pch l=0.04u w=0.8u
m22362 4512 4512 VDDPOST VDDPOST pch l=0.04u w=1u
m22363 4513 4513 VDDPOST VDDPOST pch l=0.04u w=1u
m22364 VDDREF 4480 4502 VDDREF pch l=0.04u w=0.8u
m22365 VDDREF 4481 4503 VDDREF pch l=0.04u w=0.8u
m22366 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22367 4506 4522 VDDREF VDDREF pch l=0.04u w=0.8u
m22368 4507 4523 VDDREF VDDREF pch l=0.04u w=0.8u
m22369 4508 4524 VDDREF VDDREF pch l=0.04u w=0.8u
m22370 4509 4525 VDDREF VDDREF pch l=0.04u w=0.8u
m22371 4510 4526 VDDREF VDDREF pch l=0.04u w=0.8u
m22372 VDDREF 4522 4506 VDDREF pch l=0.04u w=0.8u
m22373 VDDREF 4523 4507 VDDREF pch l=0.04u w=0.8u
m22374 VDDREF 4524 4508 VDDREF pch l=0.04u w=0.8u
m22375 VDDREF 4525 4509 VDDREF pch l=0.04u w=0.8u
m22376 VDDREF 4526 4510 VDDREF pch l=0.04u w=0.8u
m22377 VDDPOST 4515 4516 VDDPOST pch l=0.04u w=1u
m22378 VDDPOST 4518 4517 VDDPOST pch l=0.04u w=1u
m22379 4520 4502 VDDREF VDDREF pch l=0.04u w=0.8u
m22380 4521 4503 VDDREF VDDREF pch l=0.04u w=0.8u
m22381 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22382 VDDREF 4502 4520 VDDREF pch l=0.04u w=0.8u
m22383 VDDREF 4503 4521 VDDREF pch l=0.04u w=0.8u
m22384 VDDREF 4527 4522 VDDREF pch l=0.04u w=0.8u
m22385 VDDREF 4528 4523 VDDREF pch l=0.04u w=0.8u
m22386 VDDREF 4529 4524 VDDREF pch l=0.04u w=0.8u
m22387 VDDREF 4530 4525 VDDREF pch l=0.04u w=0.8u
m22388 VDDREF 4531 4526 VDDREF pch l=0.04u w=0.8u
m22389 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22390 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22391 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22392 4520 4502 VDDREF VDDREF pch l=0.04u w=0.8u
m22393 4521 4503 VDDREF VDDREF pch l=0.04u w=0.8u
m22394 VDDREF 4502 4520 VDDREF pch l=0.04u w=0.8u
m22395 VDDREF 4503 4521 VDDREF pch l=0.04u w=0.8u
m22396 4527 4497 VDDREF VDDREF pch l=0.04u w=0.8u
m22397 4528 4498 VDDREF VDDREF pch l=0.04u w=0.8u
m22398 4529 4499 VDDREF VDDREF pch l=0.04u w=0.8u
m22399 4530 4500 VDDREF VDDREF pch l=0.04u w=0.8u
m22400 4531 4501 VDDREF VDDREF pch l=0.04u w=0.8u
m22401 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22402 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22403 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22404 VDDREF 4540 4527 VDDREF pch l=0.04u w=0.8u
m22405 VDDREF 4541 4528 VDDREF pch l=0.04u w=0.8u
m22406 VDDREF 4542 4529 VDDREF pch l=0.04u w=0.8u
m22407 VDDREF 4543 4530 VDDREF pch l=0.04u w=0.8u
m22408 VDDREF 4544 4531 VDDREF pch l=0.04u w=0.8u
m22409 4532 4520 VDDREF VDDREF pch l=0.04u w=0.8u
m22410 4533 4521 VDDREF VDDREF pch l=0.04u w=0.8u
m22411 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22412 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22413 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22414 VDDREF 4520 4532 VDDREF pch l=0.04u w=0.8u
m22415 VDDREF 4521 4533 VDDREF pch l=0.04u w=0.8u
m22416 4534 4497 VDDREF VDDREF pch l=0.04u w=0.8u
m22417 4535 4498 VDDREF VDDREF pch l=0.04u w=0.8u
m22418 4536 4499 VDDREF VDDREF pch l=0.04u w=0.8u
m22419 4537 4500 VDDREF VDDREF pch l=0.04u w=0.8u
m22420 4538 4501 VDDREF VDDREF pch l=0.04u w=0.8u
m22421 4532 4520 VDDREF VDDREF pch l=0.04u w=0.8u
m22422 4533 4521 VDDREF VDDREF pch l=0.04u w=0.8u
m22423 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22424 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22425 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22426 VDDREF 4520 4532 VDDREF pch l=0.04u w=0.8u
m22427 VDDREF 4521 4533 VDDREF pch l=0.04u w=0.8u
m22428 4540 4527 VDDREF VDDREF pch l=0.04u w=0.8u
m22429 4541 4528 VDDREF VDDREF pch l=0.04u w=0.8u
m22430 4542 4529 VDDREF VDDREF pch l=0.04u w=0.8u
m22431 4543 4530 VDDREF VDDREF pch l=0.04u w=0.8u
m22432 4544 4531 VDDREF VDDREF pch l=0.04u w=0.8u
m22433 4532 4520 VDDREF VDDREF pch l=0.04u w=0.8u
m22434 4533 4521 VDDREF VDDREF pch l=0.04u w=0.8u
m22435 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22436 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22437 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22438 VDDREF 4534 4540 VDDREF pch l=0.04u w=0.8u
m22439 VDDREF 4535 4541 VDDREF pch l=0.04u w=0.8u
m22440 VDDREF 4536 4542 VDDREF pch l=0.04u w=0.8u
m22441 VDDREF 4537 4543 VDDREF pch l=0.04u w=0.8u
m22442 VDDREF 4538 4544 VDDREF pch l=0.04u w=0.8u
m22443 VDDREF 4520 4532 VDDREF pch l=0.04u w=0.8u
m22444 VDDREF 4521 4533 VDDREF pch l=0.04u w=0.8u
m22445 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22446 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22447 VDDREF 4551 VDDREF VDDREF pch l=0.26u w=1u
m22448 4545 4540 VDDREF VDDREF pch l=0.04u w=0.8u
m22449 4546 4541 VDDREF VDDREF pch l=0.04u w=0.8u
m22450 4547 4542 VDDREF VDDREF pch l=0.04u w=0.8u
m22451 4548 4543 VDDREF VDDREF pch l=0.04u w=0.8u
m22452 4549 4544 VDDREF VDDREF pch l=0.04u w=0.8u
m22453 4532 4520 VDDREF VDDREF pch l=0.04u w=0.8u
m22454 4533 4521 VDDREF VDDREF pch l=0.04u w=0.8u
m22455 4550 4550 VDDREF VDDREF pch l=0.04u w=1u
m22456 VDDREF 4520 4532 VDDREF pch l=0.04u w=0.8u
m22457 VDDREF 4521 4533 VDDREF pch l=0.04u w=0.8u
m22458 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22459 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22460 4554 4545 VDDREF VDDREF pch l=0.04u w=0.8u
m22461 4555 4546 VDDREF VDDREF pch l=0.04u w=0.8u
m22462 4556 4547 VDDREF VDDREF pch l=0.04u w=0.8u
m22463 4557 4548 VDDREF VDDREF pch l=0.04u w=0.8u
m22464 4558 4549 VDDREF VDDREF pch l=0.04u w=0.8u
m22465 4532 4520 VDDREF VDDREF pch l=0.04u w=0.8u
m22466 4533 4521 VDDREF VDDREF pch l=0.04u w=0.8u
m22467 VDDREF 4553 4552 VDDREF pch l=0.04u w=1u
m22468 VDDREF 4545 4554 VDDREF pch l=0.04u w=0.8u
m22469 VDDREF 4546 4555 VDDREF pch l=0.04u w=0.8u
m22470 VDDREF 4547 4556 VDDREF pch l=0.04u w=0.8u
m22471 VDDREF 4548 4557 VDDREF pch l=0.04u w=0.8u
m22472 VDDREF 4549 4558 VDDREF pch l=0.04u w=0.8u
m22473 VDDREF 4520 4532 VDDREF pch l=0.04u w=0.8u
m22474 VDDREF 4521 4533 VDDREF pch l=0.04u w=0.8u
m22475 VDDPOST 4559 VDDPOST VDDPOST pch l=0.26u w=1u
m22476 VDDPOST 4562 VDDPOST VDDPOST pch l=0.26u w=1u
m22477 4554 4545 VDDREF VDDREF pch l=0.04u w=0.8u
m22478 4555 4546 VDDREF VDDREF pch l=0.04u w=0.8u
m22479 4556 4547 VDDREF VDDREF pch l=0.04u w=0.8u
m22480 4557 4548 VDDREF VDDREF pch l=0.04u w=0.8u
m22481 4558 4549 VDDREF VDDREF pch l=0.04u w=0.8u
m22482 4532 4520 VDDREF VDDREF pch l=0.04u w=0.8u
m22483 4533 4521 VDDREF VDDREF pch l=0.04u w=0.8u
m22484 4560 4560 VDDPOST VDDPOST pch l=0.04u w=1u
m22485 4561 4561 VDDPOST VDDPOST pch l=0.04u w=1u
m22486 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22487 VDDREF 4545 4554 VDDREF pch l=0.04u w=0.8u
m22488 VDDREF 4546 4555 VDDREF pch l=0.04u w=0.8u
m22489 VDDREF 4547 4556 VDDREF pch l=0.04u w=0.8u
m22490 VDDREF 4548 4557 VDDREF pch l=0.04u w=0.8u
m22491 VDDREF 4549 4558 VDDREF pch l=0.04u w=0.8u
m22492 VDDREF 4520 4532 VDDREF pch l=0.04u w=0.8u
m22493 VDDREF 4521 4533 VDDREF pch l=0.04u w=0.8u
m22494 VDDPOST 4564 4565 VDDPOST pch l=0.04u w=1u
m22495 VDDPOST 4567 4566 VDDPOST pch l=0.04u w=1u
m22496 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22497 4568 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22498 4569 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22499 4570 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22500 4571 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22501 4572 4395 VDDREF VDDREF pch l=0.04u w=0.8u
m22502 4573 4606 VDDREF VDDREF pch l=0.04u w=0.8u
m22503 4574 4607 VDDREF VDDREF pch l=0.04u w=0.8u
m22504 VDDREF 2666 4568 VDDREF pch l=0.04u w=0.8u
m22505 VDDREF 2927 4569 VDDREF pch l=0.04u w=0.8u
m22506 VDDREF 3205 4570 VDDREF pch l=0.04u w=0.8u
m22507 VDDREF 4425 4571 VDDREF pch l=0.04u w=0.8u
m22508 VDDREF 3937 4572 VDDREF pch l=0.04u w=0.8u
m22509 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22510 VDDREF 4606 4573 VDDREF pch l=0.04u w=0.8u
m22511 VDDREF 4607 4574 VDDREF pch l=0.04u w=0.8u
m22512 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22513 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22514 4573 4606 VDDREF VDDREF pch l=0.04u w=0.8u
m22515 4574 4607 VDDREF VDDREF pch l=0.04u w=0.8u
m22516 4575 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22517 4576 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22518 4577 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22519 4578 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22520 4579 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22521 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22522 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22523 VDDREF 4606 4573 VDDREF pch l=0.04u w=0.8u
m22524 VDDREF 4607 4574 VDDREF pch l=0.04u w=0.8u
m22525 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22526 4573 4606 VDDREF VDDREF pch l=0.04u w=0.8u
m22527 4574 4607 VDDREF VDDREF pch l=0.04u w=0.8u
m22528 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22529 4580 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22530 4581 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22531 4582 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22532 4583 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22533 4584 DACPD VDDREF VDDREF pch l=0.04u w=0.8u
m22534 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22535 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22536 VDDREF 4606 4573 VDDREF pch l=0.04u w=0.8u
m22537 VDDREF 4607 4574 VDDREF pch l=0.04u w=0.8u
m22538 VDDREF DACPD 4580 VDDREF pch l=0.04u w=0.8u
m22539 VDDREF DACPD 4581 VDDREF pch l=0.04u w=0.8u
m22540 VDDREF DACPD 4582 VDDREF pch l=0.04u w=0.8u
m22541 VDDREF DACPD 4583 VDDREF pch l=0.04u w=0.8u
m22542 VDDREF DACPD 4584 VDDREF pch l=0.04u w=0.8u
m22543 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22544 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22545 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22546 4573 4606 VDDREF VDDREF pch l=0.04u w=0.8u
m22547 4574 4607 VDDREF VDDREF pch l=0.04u w=0.8u
m22548 4586 4575 VDDREF VDDREF pch l=0.04u w=0.8u
m22549 4587 4576 VDDREF VDDREF pch l=0.04u w=0.8u
m22550 4588 4577 VDDREF VDDREF pch l=0.04u w=0.8u
m22551 4589 4578 VDDREF VDDREF pch l=0.04u w=0.8u
m22552 4590 4579 VDDREF VDDREF pch l=0.04u w=0.8u
m22553 VDDREF 4606 4573 VDDREF pch l=0.04u w=0.8u
m22554 VDDREF 4607 4574 VDDREF pch l=0.04u w=0.8u
m22555 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22556 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22557 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22558 VDDREF 4568 4586 VDDREF pch l=0.04u w=0.8u
m22559 VDDREF 4569 4587 VDDREF pch l=0.04u w=0.8u
m22560 VDDREF 4570 4588 VDDREF pch l=0.04u w=0.8u
m22561 VDDREF 4571 4589 VDDREF pch l=0.04u w=0.8u
m22562 VDDREF 4572 4590 VDDREF pch l=0.04u w=0.8u
m22563 4573 4606 VDDREF VDDREF pch l=0.04u w=0.8u
m22564 4574 4607 VDDREF VDDREF pch l=0.04u w=0.8u
m22565 VDDREF 4606 4573 VDDREF pch l=0.04u w=0.8u
m22566 VDDREF 4607 4574 VDDREF pch l=0.04u w=0.8u
m22567 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22568 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22569 VDDREF 4597 VDDREF VDDREF pch l=0.26u w=1u
m22570 4591 4586 VDDREF VDDREF pch l=0.04u w=0.8u
m22571 4592 4587 VDDREF VDDREF pch l=0.04u w=0.8u
m22572 4593 4588 VDDREF VDDREF pch l=0.04u w=0.8u
m22573 4594 4589 VDDREF VDDREF pch l=0.04u w=0.8u
m22574 4595 4590 VDDREF VDDREF pch l=0.04u w=0.8u
m22575 4573 4606 VDDREF VDDREF pch l=0.04u w=0.8u
m22576 4574 4607 VDDREF VDDREF pch l=0.04u w=0.8u
m22577 4596 4596 VDDREF VDDREF pch l=0.04u w=1u
m22578 VDDREF 4580 4591 VDDREF pch l=0.04u w=0.8u
m22579 VDDREF 4581 4592 VDDREF pch l=0.04u w=0.8u
m22580 VDDREF 4582 4593 VDDREF pch l=0.04u w=0.8u
m22581 VDDREF 4583 4594 VDDREF pch l=0.04u w=0.8u
m22582 VDDREF 4584 4595 VDDREF pch l=0.04u w=0.8u
m22583 VDDREF 4606 4573 VDDREF pch l=0.04u w=0.8u
m22584 VDDREF 4607 4574 VDDREF pch l=0.04u w=0.8u
m22585 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22586 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22587 VDDREF 4599 4598 VDDREF pch l=0.04u w=1u
m22588 4601 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22589 4602 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22590 4603 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22591 4604 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22592 4605 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22593 4606 4624 VDDREF VDDREF pch l=0.04u w=0.8u
m22594 4607 4625 VDDREF VDDREF pch l=0.04u w=0.8u
m22595 VDDPOST 4608 VDDPOST VDDPOST pch l=0.26u w=1u
m22596 VDDPOST 4611 VDDPOST VDDPOST pch l=0.26u w=1u
m22597 VDDREF 4624 4606 VDDREF pch l=0.04u w=0.8u
m22598 VDDREF 4625 4607 VDDREF pch l=0.04u w=0.8u
m22599 4609 4609 VDDPOST VDDPOST pch l=0.04u w=1u
m22600 4610 4610 VDDPOST VDDPOST pch l=0.04u w=1u
m22601 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22602 4612 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22603 4613 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22604 4614 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22605 4615 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22606 4616 155 VDDREF VDDREF pch l=0.04u w=0.8u
m22607 4606 4624 VDDREF VDDREF pch l=0.04u w=0.8u
m22608 4607 4625 VDDREF VDDREF pch l=0.04u w=0.8u
m22609 VDDREF 4392 4612 VDDREF pch l=0.04u w=0.8u
m22610 VDDREF 4392 4613 VDDREF pch l=0.04u w=0.8u
m22611 VDDREF 4392 4614 VDDREF pch l=0.04u w=0.8u
m22612 VDDREF 4392 4615 VDDREF pch l=0.04u w=0.8u
m22613 VDDREF 4392 4616 VDDREF pch l=0.04u w=0.8u
m22614 VDDREF 4624 4606 VDDREF pch l=0.04u w=0.8u
m22615 VDDREF 4625 4607 VDDREF pch l=0.04u w=0.8u
m22616 4617 4649 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22617 FOUTVCO 4639 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22618 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22619 VDDPOST 4649 4617 VDDPOST pch l=0.04u w=0.8u
m22620 VDDPOST 4639 FOUTVCO VDDPOST pch l=0.04u w=0.8u
m22621 4619 4601 VDDREF VDDREF pch l=0.04u w=0.8u
m22622 4620 4602 VDDREF VDDREF pch l=0.04u w=0.8u
m22623 4621 4603 VDDREF VDDREF pch l=0.04u w=0.8u
m22624 4622 4604 VDDREF VDDREF pch l=0.04u w=0.8u
m22625 4623 4605 VDDREF VDDREF pch l=0.04u w=0.8u
m22626 4624 4640 VDDREF VDDREF pch l=0.04u w=0.8u
m22627 4625 4641 VDDREF VDDREF pch l=0.04u w=0.8u
m22628 4617 4649 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22629 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22630 FOUTVCO 4639 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22631 VDDREF 4591 4619 VDDREF pch l=0.04u w=0.8u
m22632 VDDREF 4592 4620 VDDREF pch l=0.04u w=0.8u
m22633 VDDREF 4593 4621 VDDREF pch l=0.04u w=0.8u
m22634 VDDREF 4594 4622 VDDREF pch l=0.04u w=0.8u
m22635 VDDREF 4595 4623 VDDREF pch l=0.04u w=0.8u
m22636 VDDREF 2426 4624 VDDREF pch l=0.04u w=0.8u
m22637 VDDREF 4426 4625 VDDREF pch l=0.04u w=0.8u
m22638 VDDPOST 4649 4617 VDDPOST pch l=0.04u w=0.8u
m22639 VDDPOST 4639 FOUTVCO VDDPOST pch l=0.04u w=0.8u
m22640 4624 2426 VDDREF VDDREF pch l=0.04u w=0.8u
m22641 4625 4426 VDDREF VDDREF pch l=0.04u w=0.8u
m22642 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22643 4617 4649 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22644 FOUTVCO 4639 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22645 VDDREF 4640 4624 VDDREF pch l=0.04u w=0.8u
m22646 VDDREF 4641 4625 VDDREF pch l=0.04u w=0.8u
m22647 4627 4619 VDDREF VDDREF pch l=0.04u w=0.8u
m22648 4628 4620 VDDREF VDDREF pch l=0.04u w=0.8u
m22649 4629 4621 VDDREF VDDREF pch l=0.04u w=0.8u
m22650 4630 4622 VDDREF VDDREF pch l=0.04u w=0.8u
m22651 4631 4623 VDDREF VDDREF pch l=0.04u w=0.8u
m22652 VDDPOST 4649 4617 VDDPOST pch l=0.04u w=0.8u
m22653 VDDPOST 4639 FOUTVCO VDDPOST pch l=0.04u w=0.8u
m22654 VDDREF 4612 4627 VDDREF pch l=0.04u w=0.8u
m22655 VDDREF 4613 4628 VDDREF pch l=0.04u w=0.8u
m22656 VDDREF 4614 4629 VDDREF pch l=0.04u w=0.8u
m22657 VDDREF 4615 4630 VDDREF pch l=0.04u w=0.8u
m22658 VDDREF 4616 4631 VDDREF pch l=0.04u w=0.8u
m22659 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22660 4617 4649 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22661 FOUTVCO 4639 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22662 4632 2426 VDDREF VDDREF pch l=0.04u w=0.8u
m22663 4633 4426 VDDREF VDDREF pch l=0.04u w=0.8u
m22664 VDDPOST 4649 4617 VDDPOST pch l=0.04u w=0.8u
m22665 VDDPOST 4639 FOUTVCO VDDPOST pch l=0.04u w=0.8u
m22666 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22667 4634 4627 VDDREF VDDREF pch l=0.04u w=0.8u
m22668 4635 4628 VDDREF VDDREF pch l=0.04u w=0.8u
m22669 4636 4629 VDDREF VDDREF pch l=0.04u w=0.8u
m22670 4637 4630 VDDREF VDDREF pch l=0.04u w=0.8u
m22671 4638 4631 VDDREF VDDREF pch l=0.04u w=0.8u
m22672 4640 4624 VDDREF VDDREF pch l=0.04u w=0.8u
m22673 4641 4625 VDDREF VDDREF pch l=0.04u w=0.8u
m22674 4642 4649 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22675 VDDPOST 4642 4639 VDDPOST pch l=0.04u w=0.8u
m22676 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22677 VDDREF 4632 4640 VDDREF pch l=0.04u w=0.8u
m22678 VDDREF 4633 4641 VDDREF pch l=0.04u w=0.8u
m22679 4644 4659 VDDREF VDDREF pch l=0.04u w=0.8u
m22680 4645 4660 VDDREF VDDREF pch l=0.04u w=0.8u
m22681 4646 4661 VDDREF VDDREF pch l=0.04u w=0.8u
m22682 4647 4662 VDDREF VDDREF pch l=0.04u w=0.8u
m22683 4648 4663 VDDREF VDDREF pch l=0.04u w=0.8u
m22684 VDDPOST 4649 4642 VDDPOST pch l=0.04u w=0.8u
m22685 4639 4642 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22686 4640 4632 VDDREF VDDREF pch l=0.04u w=0.8u
m22687 4641 4633 VDDREF VDDREF pch l=0.04u w=0.8u
m22688 VDDREF 4659 4644 VDDREF pch l=0.04u w=0.8u
m22689 VDDREF 4660 4645 VDDREF pch l=0.04u w=0.8u
m22690 VDDREF 4661 4646 VDDREF pch l=0.04u w=0.8u
m22691 VDDREF 4662 4647 VDDREF pch l=0.04u w=0.8u
m22692 VDDREF 4663 4648 VDDREF pch l=0.04u w=0.8u
m22693 VDDPOST 4687 4639 VDDPOST pch l=0.04u w=0.8u
m22694 VDDREF 4652 VDDREF VDDREF pch l=0.26u w=1u
m22695 VDDREF 4624 4640 VDDREF pch l=0.04u w=0.8u
m22696 VDDREF 4625 4641 VDDREF pch l=0.04u w=0.8u
m22697 4644 4659 VDDREF VDDREF pch l=0.04u w=0.8u
m22698 4645 4660 VDDREF VDDREF pch l=0.04u w=0.8u
m22699 4646 4661 VDDREF VDDREF pch l=0.04u w=0.8u
m22700 4647 4662 VDDREF VDDREF pch l=0.04u w=0.8u
m22701 4648 4663 VDDREF VDDREF pch l=0.04u w=0.8u
m22702 4649 4679 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22703 4651 4651 VDDREF VDDREF pch l=0.04u w=1u
m22704 VDDREF 4659 4644 VDDREF pch l=0.04u w=0.8u
m22705 VDDREF 4660 4645 VDDREF pch l=0.04u w=0.8u
m22706 VDDREF 4661 4646 VDDREF pch l=0.04u w=0.8u
m22707 VDDREF 4662 4647 VDDREF pch l=0.04u w=0.8u
m22708 VDDREF 4663 4648 VDDREF pch l=0.04u w=0.8u
m22709 VDDPOST 4679 4649 VDDPOST pch l=0.04u w=0.8u
m22710 4654 4699 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22711 4657 4640 VDDREF VDDREF pch l=0.04u w=0.8u
m22712 4658 4641 VDDREF VDDREF pch l=0.04u w=0.8u
m22713 4649 4679 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22714 VDDPOST 4642 4654 VDDPOST pch l=0.04u w=0.8u
m22715 VDDREF 4656 4655 VDDREF pch l=0.04u w=1u
m22716 VDDREF 4640 4657 VDDREF pch l=0.04u w=0.8u
m22717 VDDREF 4641 4658 VDDREF pch l=0.04u w=0.8u
m22718 VDDREF 4664 4659 VDDREF pch l=0.04u w=0.8u
m22719 VDDREF 4665 4660 VDDREF pch l=0.04u w=0.8u
m22720 VDDREF 4666 4661 VDDREF pch l=0.04u w=0.8u
m22721 VDDREF 4667 4662 VDDREF pch l=0.04u w=0.8u
m22722 VDDREF 4668 4663 VDDREF pch l=0.04u w=0.8u
m22723 VDDPOST 4679 4649 VDDPOST pch l=0.04u w=0.8u
m22724 4654 4642 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22725 4657 4640 VDDREF VDDREF pch l=0.04u w=0.8u
m22726 4658 4641 VDDREF VDDREF pch l=0.04u w=0.8u
m22727 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22728 VDDREF 4640 4657 VDDREF pch l=0.04u w=0.8u
m22729 VDDREF 4641 4658 VDDREF pch l=0.04u w=0.8u
m22730 4664 4634 VDDREF VDDREF pch l=0.04u w=0.8u
m22731 4665 4635 VDDREF VDDREF pch l=0.04u w=0.8u
m22732 4666 4636 VDDREF VDDREF pch l=0.04u w=0.8u
m22733 4667 4637 VDDREF VDDREF pch l=0.04u w=0.8u
m22734 4668 4638 VDDREF VDDREF pch l=0.04u w=0.8u
m22735 4669 4654 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22736 VDDREF 4682 4664 VDDREF pch l=0.04u w=0.8u
m22737 VDDREF 4683 4665 VDDREF pch l=0.04u w=0.8u
m22738 VDDREF 4684 4666 VDDREF pch l=0.04u w=0.8u
m22739 VDDREF 4685 4667 VDDREF pch l=0.04u w=0.8u
m22740 VDDREF 4686 4668 VDDREF pch l=0.04u w=0.8u
m22741 VDDPOST 4654 4669 VDDPOST pch l=0.04u w=0.8u
m22742 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22743 4671 4657 VDDREF VDDREF pch l=0.04u w=0.8u
m22744 4672 4658 VDDREF VDDREF pch l=0.04u w=0.8u
m22745 4669 4654 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22746 VDDREF 4657 4671 VDDREF pch l=0.04u w=0.8u
m22747 VDDREF 4658 4672 VDDREF pch l=0.04u w=0.8u
m22748 4679 4680 36642 VDDPOST pch l=0.225u w=0.15u
m22749 VDDPOST 4680 36642 VDDPOST pch l=0.225u w=0.15u
m22750 4674 4634 VDDREF VDDREF pch l=0.04u w=0.8u
m22751 4675 4635 VDDREF VDDREF pch l=0.04u w=0.8u
m22752 4676 4636 VDDREF VDDREF pch l=0.04u w=0.8u
m22753 4677 4637 VDDREF VDDREF pch l=0.04u w=0.8u
m22754 4678 4638 VDDREF VDDREF pch l=0.04u w=0.8u
m22755 VDDPOST 4654 4669 VDDPOST pch l=0.04u w=0.8u
m22756 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22757 4671 4657 VDDREF VDDREF pch l=0.04u w=0.8u
m22758 4672 4658 VDDREF VDDREF pch l=0.04u w=0.8u
m22759 4669 4654 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22760 VDDREF 4657 4671 VDDREF pch l=0.04u w=0.8u
m22761 VDDREF 4658 4672 VDDREF pch l=0.04u w=0.8u
m22762 VDDPOST 4654 4669 VDDPOST pch l=0.04u w=0.8u
m22763 4682 4664 VDDREF VDDREF pch l=0.04u w=0.8u
m22764 4683 4665 VDDREF VDDREF pch l=0.04u w=0.8u
m22765 4684 4666 VDDREF VDDREF pch l=0.04u w=0.8u
m22766 4685 4667 VDDREF VDDREF pch l=0.04u w=0.8u
m22767 4686 4668 VDDREF VDDREF pch l=0.04u w=0.8u
m22768 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22769 4671 4657 VDDREF VDDREF pch l=0.04u w=0.8u
m22770 4672 4658 VDDREF VDDREF pch l=0.04u w=0.8u
m22771 4669 4654 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22772 VDDREF 4674 4682 VDDREF pch l=0.04u w=0.8u
m22773 VDDREF 4675 4683 VDDREF pch l=0.04u w=0.8u
m22774 VDDREF 4676 4684 VDDREF pch l=0.04u w=0.8u
m22775 VDDREF 4677 4685 VDDREF pch l=0.04u w=0.8u
m22776 VDDREF 4678 4686 VDDREF pch l=0.04u w=0.8u
m22777 VDDPOST 4693 4679 VDDPOST pch l=0.04u w=0.8u
m22778 VDDREF 4657 4671 VDDREF pch l=0.04u w=0.8u
m22779 VDDREF 4658 4672 VDDREF pch l=0.04u w=0.8u
m22780 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22781 VDDPOST 4654 4669 VDDPOST pch l=0.04u w=0.8u
m22782 4679 4693 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22783 VDDPOST 4693 4679 VDDPOST pch l=0.04u w=0.8u
m22784 4688 4682 VDDREF VDDREF pch l=0.04u w=0.8u
m22785 4689 4683 VDDREF VDDREF pch l=0.04u w=0.8u
m22786 4690 4684 VDDREF VDDREF pch l=0.04u w=0.8u
m22787 4691 4685 VDDREF VDDREF pch l=0.04u w=0.8u
m22788 4692 4686 VDDREF VDDREF pch l=0.04u w=0.8u
m22789 4671 4657 VDDREF VDDREF pch l=0.04u w=0.8u
m22790 4672 4658 VDDREF VDDREF pch l=0.04u w=0.8u
m22791 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22792 37078 FOUTVCOPD 4687 VDDPOST pch l=0.04u w=0.8u
m22793 VDDREF 4657 4671 VDDREF pch l=0.04u w=0.8u
m22794 VDDREF 4658 4672 VDDREF pch l=0.04u w=0.8u
m22795 VDDPOST PD 37078 VDDPOST pch l=0.04u w=0.8u
m22796 VDDPOST 4693 4693 VDDPOST pch l=0.04u w=0.65u
m22797 4694 4688 VDDREF VDDREF pch l=0.04u w=0.8u
m22798 4695 4689 VDDREF VDDREF pch l=0.04u w=0.8u
m22799 4696 4690 VDDREF VDDREF pch l=0.04u w=0.8u
m22800 4697 4691 VDDREF VDDREF pch l=0.04u w=0.8u
m22801 4698 4692 VDDREF VDDREF pch l=0.04u w=0.8u
m22802 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22803 4671 4657 VDDREF VDDREF pch l=0.04u w=0.8u
m22804 4672 4658 VDDREF VDDREF pch l=0.04u w=0.8u
m22805 VDDREF 4688 4694 VDDREF pch l=0.04u w=0.8u
m22806 VDDREF 4689 4695 VDDREF pch l=0.04u w=0.8u
m22807 VDDREF 4690 4696 VDDREF pch l=0.04u w=0.8u
m22808 VDDREF 4691 4697 VDDREF pch l=0.04u w=0.8u
m22809 VDDREF 4692 4698 VDDREF pch l=0.04u w=0.8u
m22810 VDDREF 4657 4671 VDDREF pch l=0.04u w=0.8u
m22811 VDDREF 4658 4672 VDDREF pch l=0.04u w=0.8u
m22812 37439 PD VDDPOST VDDPOST pch l=0.04u w=0.8u
m22813 4694 4688 VDDREF VDDREF pch l=0.04u w=0.8u
m22814 4695 4689 VDDREF VDDREF pch l=0.04u w=0.8u
m22815 4696 4690 VDDREF VDDREF pch l=0.04u w=0.8u
m22816 4697 4691 VDDREF VDDREF pch l=0.04u w=0.8u
m22817 4698 4692 VDDREF VDDREF pch l=0.04u w=0.8u
m22818 VDDREF 4702 VDDREF VDDREF pch l=0.26u w=1u
m22819 4671 4657 VDDREF VDDREF pch l=0.04u w=0.8u
m22820 4672 4658 VDDREF VDDREF pch l=0.04u w=0.8u
m22821 4699 FOUTPOSTDIVPD 37439 VDDPOST pch l=0.04u w=0.8u
m22822 VDDREF 4688 4694 VDDREF pch l=0.04u w=0.8u
m22823 VDDREF 4689 4695 VDDREF pch l=0.04u w=0.8u
m22824 VDDREF 4690 4696 VDDREF pch l=0.04u w=0.8u
m22825 VDDREF 4691 4697 VDDREF pch l=0.04u w=0.8u
m22826 VDDREF 4692 4698 VDDREF pch l=0.04u w=0.8u
m22827 4701 4701 VDDREF VDDREF pch l=0.04u w=1u
m22828 VDDREF 4657 4671 VDDREF pch l=0.04u w=0.8u
m22829 VDDREF 4658 4672 VDDREF pch l=0.04u w=0.8u
m22830 4703 FOUTPOSTDIVPD VDDPOST VDDPOST pch l=0.04u w=0.8u
m22831 4704 4703 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22832 4705 4669 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22833 VDDPOST 12 4704 VDDPOST pch l=0.04u w=0.8u
m22834 VDDPOST 4669 4705 VDDPOST pch l=0.04u w=0.8u
m22835 4673 4670 4 4 pch l=0.04u w=0.8u
m22836 4707 4704 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22837 4 4670 4673 4 pch l=0.04u w=0.8u
m22838 VDDPOST 4704 4707 VDDPOST pch l=0.04u w=0.8u
m22839 4708 4788 VDDPOST VDDPOST pch l=0.04u w=0.4u
m22840 4670 4929 4 4 pch l=0.04u w=0.8u
m22841 VDDPOST 4669 4708 VDDPOST pch l=0.04u w=0.4u
m22842 40127 POSTDIV2[1] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22843 4 4929 4670 4 pch l=0.04u w=0.8u
m22844 4708 4669 VDDPOST VDDPOST pch l=0.04u w=0.4u
m22845 4709 POSTDIV2[2] 40127 VDDPOST pch l=0.04u w=0.8u
m22846 VDDPOST 4669 4708 VDDPOST pch l=0.04u w=0.4u
m22847 4708 4669 VDDPOST VDDPOST pch l=0.04u w=0.4u
m22848 4710 4709 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22849 VDDPOST 4669 4708 VDDPOST pch l=0.04u w=0.4u
m22850 4708 4669 VDDPOST VDDPOST pch l=0.04u w=0.4u
m22851 40819 4860 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22852 4 4 4 4 pch l=0.2u w=1.5u
m22853 VDDPOST 4669 4708 VDDPOST pch l=0.04u w=0.4u
m22854 4711 4710 40819 VDDPOST pch l=0.04u w=0.8u
m22855 4712 4929 4 4 pch l=0.2u w=1.5u
m22856 4708 4669 VDDPOST VDDPOST pch l=0.04u w=0.4u
m22857 4713 4953 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22858 4714 POSTDIV2[0] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22859 4 4929 4712 4 pch l=0.2u w=1.5u
m22860 41225 POSTDIV1[1] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22861 VDDPOST POSTDIV2[1] 4714 VDDPOST pch l=0.04u w=0.8u
m22862 4712 4929 4 4 pch l=0.2u w=1.5u
m22863 4715 POSTDIV1[2] 41225 VDDPOST pch l=0.04u w=0.8u
m22864 VDDPOST 4787 4716 VDDPOST pch l=0.04u w=0.8u
m22865 41399 POSTDIV2[0] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22866 4 4929 4712 4 pch l=0.2u w=1.5u
m22867 4788 4709 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22868 4786 POSTDIV2[1] 41399 VDDPOST pch l=0.04u w=0.8u
m22869 4787 4790 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22870 VDDPOST 4715 4788 VDDPOST pch l=0.04u w=0.8u
m22871 4712 4929 4 4 pch l=0.2u w=1.5u
m22872 VDDPOST 4713 4787 VDDPOST pch l=0.04u w=0.8u
m22873 4789 POSTDIV2[2] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22874 4 4929 4712 4 pch l=0.2u w=1.5u
m22875 41613 4860 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22876 VDDPOST 4793 4790 VDDPOST pch l=0.04u w=0.8u
m22877 4791 4788 41613 VDDPOST pch l=0.04u w=0.8u
m22878 4712 4929 4 4 pch l=0.2u w=1.5u
m22879 41658 4789 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22880 41675 4716 VDDPOST VDDPOST pch l=0.04u w=0.24u
m22881 4792 4714 41658 VDDPOST pch l=0.04u w=0.8u
m22882 4 4929 4712 4 pch l=0.2u w=1.5u
m22883 4793 4981 41675 VDDPOST pch l=0.04u w=0.24u
m22884 41710 BYPASS VDDPOST VDDPOST pch l=0.04u w=0.8u
m22885 4857 4874 4793 VDDPOST pch l=0.04u w=0.8u
m22886 4794 FOUTPOSTDIVPD 41710 VDDPOST pch l=0.04u w=0.8u
m22887 4712 4929 4 4 pch l=0.2u w=1.5u
m22888 4858 4789 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22889 VDDPOST 4714 4858 VDDPOST pch l=0.04u w=0.8u
m22890 4 4929 4712 4 pch l=0.2u w=1.5u
m22891 4857 4870 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22892 4860 4794 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22893 VDDPOST 4713 4857 VDDPOST pch l=0.04u w=0.8u
m22894 41953 4789 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22895 4712 4929 4 4 pch l=0.2u w=1.5u
m22896 41970 4857 VDDPOST VDDPOST pch l=0.04u w=0.12u
m22897 4866 POSTDIV1[0] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22898 4863 4786 41953 VDDPOST pch l=0.04u w=0.8u
m22899 4870 4874 41970 VDDPOST pch l=0.04u w=0.12u
m22900 4 4929 4712 4 pch l=0.2u w=1.5u
m22901 4871 4981 4870 VDDPOST pch l=0.04u w=0.8u
m22902 4872 POSTDIV1[1] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22903 4873 POSTDIV2[1] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22904 4712 4929 4 4 pch l=0.2u w=1.5u
m22905 4874 4981 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22906 4 4929 4712 4 pch l=0.2u w=1.5u
m22907 4875 POSTDIV1[2] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22908 42233 POSTDIV2[0] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22909 42269 4873 42233 VDDPOST pch l=0.04u w=0.8u
m22910 4712 4929 4 4 pch l=0.2u w=1.5u
m22911 VDDPOST 4926 4871 VDDPOST pch l=0.04u w=0.8u
m22912 42307 POSTDIV1[0] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22913 4876 4789 42269 VDDPOST pch l=0.04u w=0.8u
m22914 4 4929 4712 4 pch l=0.2u w=1.5u
m22915 42346 4872 42307 VDDPOST pch l=0.04u w=0.8u
m22916 4925 POSTDIV1[2] 42346 VDDPOST pch l=0.04u w=0.8u
m22917 4926 4931 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22918 4928 4792 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22919 4929 4974 4 4 pch l=0.2u w=1.5u
m22920 VDDPOST 4713 4926 VDDPOST pch l=0.04u w=0.8u
m22921 VDDPOST 5527 4928 VDDPOST pch l=0.04u w=0.8u
m22922 4 4974 4929 4 pch l=0.2u w=1.5u
m22923 4930 4866 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22924 4928 5527 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22925 VDDPOST 4872 4930 VDDPOST pch l=0.04u w=0.8u
m22926 VDDPOST 4934 4931 VDDPOST pch l=0.04u w=0.8u
m22927 4929 4974 4 4 pch l=0.2u w=1.5u
m22928 4930 POSTDIV1[2] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22929 42531 4871 VDDPOST VDDPOST pch l=0.04u w=0.24u
m22930 4932 4928 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22931 4934 4981 42531 VDDPOST pch l=0.04u w=0.24u
m22932 4 4974 4929 4 pch l=0.2u w=1.5u
m22933 4936 4951 4934 VDDPOST pch l=0.04u w=0.8u
m22934 4933 4930 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22935 4937 4928 4935 VDDPOST pch l=0.04u w=0.8u
m22936 4929 4974 4 4 pch l=0.2u w=1.5u
m22937 4939 4939 VDDREF VDDREF pch l=0.04u w=1u
m22938 VDDPOST 4941 4933 VDDPOST pch l=0.04u w=0.8u
m22939 43012 4932 4937 VDDPOST pch l=0.04u w=0.12u
m22940 4936 4945 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22941 4 4974 4929 4 pch l=0.2u w=1.5u
m22942 VDDPOST 4942 43012 VDDPOST pch l=0.04u w=0.12u
m22943 VDDREF PD 4940 VDDREF pch l=0.04u w=0.8u
m22944 VDDPOST 4713 4936 VDDPOST pch l=0.04u w=0.8u
m22945 4941 POSTDIV1[0] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22946 4942 4937 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22947 4943 4940 VDDREF VDDREF pch l=0.04u w=0.8u
m22948 4929 4974 4 4 pch l=0.2u w=1.5u
m22949 43379 4936 VDDPOST VDDPOST pch l=0.04u w=0.12u
m22950 VDDPOST POSTDIV1[1] 4941 VDDPOST pch l=0.04u w=0.8u
m22951 43470 FOUT4PHASEPD VDDPOST VDDPOST pch l=0.04u w=0.8u
m22952 4945 4951 43379 VDDPOST pch l=0.04u w=0.12u
m22953 4941 4875 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22954 4 4974 4929 4 pch l=0.2u w=1.5u
m22955 4947 4932 4942 VDDPOST pch l=0.04u w=0.8u
m22956 43616 FOUTPOSTDIVPD 43470 VDDPOST pch l=0.04u w=0.8u
m22957 4713 4981 4945 VDDPOST pch l=0.04u w=0.8u
m22958 43667 4928 4947 VDDPOST pch l=0.04u w=0.12u
m22959 4944 PD 43616 VDDPOST pch l=0.04u w=0.8u
m22960 4929 4974 4 4 pch l=0.2u w=1.5u
m22961 4950 POSTDIV1[0] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22962 VDDPOST 4952 43667 VDDPOST pch l=0.04u w=0.12u
m22963 4951 4981 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22964 VDDPOST 4872 4950 VDDPOST pch l=0.04u w=0.8u
m22965 4952 4947 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22966 4 4974 4929 4 pch l=0.2u w=1.5u
m22967 4953 4944 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22968 4950 POSTDIV1[2] VDDPOST VDDPOST pch l=0.04u w=0.8u
m22969 4929 4974 4 4 pch l=0.2u w=1.5u
m22970 FOUT1PH270 4970 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22971 4958 4958 VDDREF VDDREF pch l=0.04u w=1u
m22972 4959 4953 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22973 4960 4792 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22974 VDDPOST 4970 FOUT1PH270 VDDPOST pch l=0.04u w=0.8u
m22975 4956 4950 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22976 4 4974 4929 4 pch l=0.2u w=1.5u
m22977 FOUT1PH270 4970 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22978 VDDPOST 4968 4956 VDDPOST pch l=0.04u w=0.8u
m22979 VDDREF 1580 4961 VDDREF pch l=0.04u w=0.8u
m22980 4963 4792 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22981 VDDPOST 4970 FOUT1PH270 VDDPOST pch l=0.04u w=0.8u
m22982 4929 4974 4 4 pch l=0.2u w=1.5u
m22983 4964 4961 VDDREF VDDREF pch l=0.04u w=0.8u
m22984 VDDPOST 4966 4962 VDDPOST pch l=0.04u w=0.8u
m22985 VDDPOST 4952 4963 VDDPOST pch l=0.04u w=0.8u
m22986 FOUT1PH270 4970 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22987 4965 4968 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22988 4 4974 4929 4 pch l=0.2u w=1.5u
m22989 VDDPOST 4970 FOUT1PH270 VDDPOST pch l=0.04u w=0.8u
m22990 4966 4969 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22991 4967 4960 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22992 FOUT1PH270 4970 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22993 4968 4866 VDDPOST VDDPOST pch l=0.04u w=0.8u
m22994 4929 4974 4 4 pch l=0.2u w=1.5u
m22995 VDDPOST 4959 4966 VDDPOST pch l=0.04u w=0.8u
m22996 VDDPOST 4935 4967 VDDPOST pch l=0.04u w=0.8u
m22997 VDDPOST 4970 FOUT1PH270 VDDPOST pch l=0.04u w=0.8u
m22998 VDDPOST POSTDIV1[1] 4968 VDDPOST pch l=0.04u w=0.8u
m22999 4 4974 4929 4 pch l=0.2u w=1.5u
m23000 4968 POSTDIV1[2] VDDPOST VDDPOST pch l=0.04u w=0.8u
m23001 VDDPOST 4978 4969 VDDPOST pch l=0.04u w=0.8u
m23002 4972 4967 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23003 VDDPOST 5424 4970 VDDPOST pch l=0.04u w=0.8u
m23004 4974 4712 4 4 pch l=0.2u w=1.5u
m23005 45495 4962 VDDPOST VDDPOST pch l=0.04u w=0.24u
m23006 VDDPOST 4963 4972 VDDPOST pch l=0.04u w=0.8u
m23007 4970 5424 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23008 4976 4976 VDDREF VDDREF pch l=0.04u w=1u
m23009 45544 4866 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23010 4978 5143 45495 VDDPOST pch l=0.04u w=0.24u
m23011 4 4712 4974 4 pch l=0.2u w=1.5u
m23012 4972 4963 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23013 VDDPOST 4716 4970 VDDPOST pch l=0.04u w=0.8u
m23014 45696 4872 45544 VDDPOST pch l=0.04u w=0.8u
m23015 4980 4997 4978 VDDPOST pch l=0.04u w=0.8u
m23016 VDDPOST 4967 4972 VDDPOST pch l=0.04u w=0.8u
m23017 VDDREF 1487 4979 VDDREF pch l=0.04u w=0.8u
m23018 4977 4875 45696 VDDPOST pch l=0.04u w=0.8u
m23019 4974 4712 4 4 pch l=0.2u w=1.5u
m23020 VDDPOST 4986 4981 VDDPOST pch l=0.04u w=0.8u
m23021 4983 4979 VDDREF VDDREF pch l=0.04u w=0.8u
m23022 4980 4990 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23023 4985 4863 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23024 4986 5424 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23025 4 4712 4974 4 pch l=0.2u w=1.5u
m23026 VDDPOST 4959 4980 VDDPOST pch l=0.04u w=0.8u
m23027 VDDPOST 5527 4985 VDDPOST pch l=0.04u w=0.8u
m23028 4974 4712 4 4 pch l=0.2u w=1.5u
m23029 46657 4980 VDDPOST VDDPOST pch l=0.04u w=0.12u
m23030 4985 5527 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23031 4987 FOUT1PH270 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23032 4989 4977 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23033 4990 4997 46657 VDDPOST pch l=0.04u w=0.12u
m23034 VDDPOST FOUT1PH270 4987 VDDPOST pch l=0.04u w=0.8u
m23035 4 4712 4974 4 pch l=0.2u w=1.5u
m23036 VDDPOST 4708 4989 VDDPOST pch l=0.04u w=0.4u
m23037 4993 5143 4990 VDDPOST pch l=0.04u w=0.8u
m23038 4987 FOUT1PH270 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23039 4989 4708 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23040 4995 4985 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23041 4974 4712 4 4 pch l=0.2u w=1.5u
m23042 VDDPOST FOUT1PH270 4987 VDDPOST pch l=0.04u w=0.8u
m23043 VDDPOST 4708 4989 VDDPOST pch l=0.04u w=0.4u
m23044 4997 5143 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23045 4989 4708 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23046 4 4712 4974 4 pch l=0.2u w=1.5u
m23047 4998 4985 4972 VDDPOST pch l=0.04u w=0.8u
m23048 4999 4953 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23049 VDDPOST 4708 4989 VDDPOST pch l=0.04u w=0.4u
m23050 47301 4995 4998 VDDPOST pch l=0.04u w=0.12u
m23051 4974 4712 4 4 pch l=0.2u w=1.5u
m23052 4989 4708 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23053 VDDPOST 5018 4993 VDDPOST pch l=0.04u w=0.8u
m23054 VDDPOST 5019 47301 VDDPOST pch l=0.04u w=0.12u
m23055 5002 4432 5015 5014 pch l=0.04u w=0.4u
m23056 5003 4432 4 5014 pch l=0.04u w=0.4u
m23057 5004 4432 5015 5014 pch l=0.04u w=0.4u
m23058 5005 4432 4 5014 pch l=0.04u w=0.4u
m23059 5006 4432 5015 5014 pch l=0.04u w=0.4u
m23060 5007 4432 4 5014 pch l=0.04u w=0.4u
m23061 5008 4432 5015 5014 pch l=0.04u w=0.4u
m23062 5009 4432 4 5014 pch l=0.04u w=0.4u
m23063 5010 4432 5015 5014 pch l=0.04u w=0.4u
m23064 5011 4432 4 5014 pch l=0.04u w=0.4u
m23065 5012 4433 4 5014 pch l=0.04u w=0.4u
m23066 5013 4433 4 5014 pch l=0.04u w=0.4u
m23067 VDDPOST 4708 4989 VDDPOST pch l=0.04u w=0.4u
m23068 5019 4998 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23069 4 4712 4974 4 pch l=0.2u w=1.5u
m23070 VSS 4532 5002 5014 pch l=0.04u w=0.4u
m23071 5015 4532 5003 5014 pch l=0.04u w=0.4u
m23072 VSS 4532 5004 5014 pch l=0.04u w=0.4u
m23073 5015 4532 5005 5014 pch l=0.04u w=0.4u
m23074 VSS 4532 5006 5014 pch l=0.04u w=0.4u
m23075 5015 4532 5007 5014 pch l=0.04u w=0.4u
m23076 VSS 4532 5008 5014 pch l=0.04u w=0.4u
m23077 5015 4532 5009 5014 pch l=0.04u w=0.4u
m23078 VSS 4532 5010 5014 pch l=0.04u w=0.4u
m23079 5015 4532 5011 5014 pch l=0.04u w=0.4u
m23080 5015 4533 5012 5014 pch l=0.04u w=0.4u
m23081 5015 4533 5013 5014 pch l=0.04u w=0.4u
m23082 4989 4708 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23083 VDDPOST 5021 5017 VDDPOST pch l=0.04u w=0.8u
m23084 5018 5023 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23085 4974 4712 4 4 pch l=0.2u w=1.5u
m23086 VDDPOST 4959 5018 VDDPOST pch l=0.04u w=0.8u
m23087 5022 4995 5019 VDDPOST pch l=0.04u w=0.8u
m23088 5021 5039 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23089 VDDREF 5037 5016 VDDREF pch l=0.26u w=0.4u
m23090 5024 4989 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23091 47686 4985 5022 VDDPOST pch l=0.04u w=0.12u
m23092 4 4712 4974 4 pch l=0.2u w=1.5u
m23093 VDDPOST 4999 5021 VDDPOST pch l=0.04u w=0.8u
m23094 VDDPOST 5045 5023 VDDPOST pch l=0.04u w=0.8u
m23095 VDDPOST 5042 47686 VDDPOST pch l=0.04u w=0.12u
m23096 4974 4712 4 4 pch l=0.2u w=1.5u
m23097 5025 4671 5015 5014 pch l=0.04u w=0.4u
m23098 5026 4671 4 5014 pch l=0.04u w=0.4u
m23099 5027 4671 5015 5014 pch l=0.04u w=0.4u
m23100 5028 4671 4 5014 pch l=0.04u w=0.4u
m23101 5029 4671 5015 5014 pch l=0.04u w=0.4u
m23102 5030 4671 4 5014 pch l=0.04u w=0.4u
m23103 5031 4671 5015 5014 pch l=0.04u w=0.4u
m23104 5032 4671 4 5014 pch l=0.04u w=0.4u
m23105 5033 4671 5015 5014 pch l=0.04u w=0.4u
m23106 5034 4671 4 5014 pch l=0.04u w=0.4u
m23107 5035 4672 4 5014 pch l=0.04u w=0.4u
m23108 5036 4672 4 5014 pch l=0.04u w=0.4u
m23109 47861 4993 VDDPOST VDDPOST pch l=0.04u w=0.24u
m23110 VDDREF 2426 5037 VDDREF pch l=0.04u w=0.8u
m23111 5042 5022 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23112 5041 4989 5038 VDDPOST pch l=0.04u w=0.8u
m23113 VSS 4573 5025 5014 pch l=0.04u w=0.4u
m23114 5015 4573 5026 5014 pch l=0.04u w=0.4u
m23115 VSS 4573 5027 5014 pch l=0.04u w=0.4u
m23116 5015 4573 5028 5014 pch l=0.04u w=0.4u
m23117 VSS 4573 5029 5014 pch l=0.04u w=0.4u
m23118 5015 4573 5030 5014 pch l=0.04u w=0.4u
m23119 VSS 4573 5031 5014 pch l=0.04u w=0.4u
m23120 5015 4573 5032 5014 pch l=0.04u w=0.4u
m23121 VSS 4573 5033 5014 pch l=0.04u w=0.4u
m23122 5015 4573 5034 5014 pch l=0.04u w=0.4u
m23123 5015 4574 5035 5014 pch l=0.04u w=0.4u
m23124 5015 4574 5036 5014 pch l=0.04u w=0.4u
m23125 5045 5143 47861 VDDPOST pch l=0.04u w=0.24u
m23126 VDDPOST 5049 5039 VDDPOST pch l=0.04u w=0.8u
m23127 5044 5037 VDDREF VDDREF pch l=0.04u w=0.8u
m23128 47931 5024 5041 VDDPOST pch l=0.04u w=0.12u
m23129 4 4712 4974 4 pch l=0.2u w=1.5u
m23130 5046 5088 5045 VDDPOST pch l=0.04u w=0.8u
m23131 47986 5017 VDDPOST VDDPOST pch l=0.04u w=0.24u
m23132 VDDPOST 5051 47931 VDDPOST pch l=0.04u w=0.12u
m23133 5047 4863 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23134 4974 4712 4 4 pch l=0.2u w=1.5u
m23135 5049 5248 47986 VDDPOST pch l=0.04u w=0.24u
m23136 5051 5041 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23137 5064 5094 5049 VDDPOST pch l=0.04u w=0.8u
m23138 5050 5044 VDDREF VDDREF pch l=0.26u w=0.4u
m23139 5046 5069 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23140 4 4712 4974 4 pch l=0.2u w=1.5u
m23141 5065 4863 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23142 5052 4432 5015 5014 pch l=0.04u w=0.4u
m23143 5053 4432 4 5014 pch l=0.04u w=0.4u
m23144 5054 4432 5015 5014 pch l=0.04u w=0.4u
m23145 5055 4432 4 5014 pch l=0.04u w=0.4u
m23146 5056 4432 5015 5014 pch l=0.04u w=0.4u
m23147 5057 4432 4 5014 pch l=0.04u w=0.4u
m23148 5058 4432 5015 5014 pch l=0.04u w=0.4u
m23149 5059 4432 4 5014 pch l=0.04u w=0.4u
m23150 5060 4432 5015 5014 pch l=0.04u w=0.4u
m23151 5061 4432 4 5014 pch l=0.04u w=0.4u
m23152 5062 4433 4 5014 pch l=0.04u w=0.4u
m23153 5063 4433 4 5014 pch l=0.04u w=0.4u
m23154 VDDPOST 4959 5046 VDDPOST pch l=0.04u w=0.8u
m23155 5066 5024 5051 VDDPOST pch l=0.04u w=0.8u
m23156 VDDPOST 5042 5065 VDDPOST pch l=0.04u w=0.8u
m23157 VSS 4532 5052 5014 pch l=0.04u w=0.4u
m23158 5015 4532 5053 5014 pch l=0.04u w=0.4u
m23159 VSS 4532 5054 5014 pch l=0.04u w=0.4u
m23160 5015 4532 5055 5014 pch l=0.04u w=0.4u
m23161 VSS 4532 5056 5014 pch l=0.04u w=0.4u
m23162 5015 4532 5057 5014 pch l=0.04u w=0.4u
m23163 VSS 4532 5058 5014 pch l=0.04u w=0.4u
m23164 5015 4532 5059 5014 pch l=0.04u w=0.4u
m23165 VSS 4532 5060 5014 pch l=0.04u w=0.4u
m23166 5015 4532 5061 5014 pch l=0.04u w=0.4u
m23167 5015 4533 5062 5014 pch l=0.04u w=0.4u
m23168 5015 4533 5063 5014 pch l=0.04u w=0.4u
m23169 48288 5046 VDDPOST VDDPOST pch l=0.04u w=0.12u
m23170 5064 5085 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23171 4 4 4 4 pch l=0.2u w=1.5u
m23172 48327 4989 5066 VDDPOST pch l=0.04u w=0.12u
m23173 5069 5088 48288 VDDPOST pch l=0.04u w=0.12u
m23174 VDDPOST 4999 5064 VDDPOST pch l=0.04u w=0.8u
m23175 VDDPOST 5071 48327 VDDPOST pch l=0.04u w=0.12u
m23176 5070 5047 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23177 4959 5143 5069 VDDPOST pch l=0.04u w=0.8u
m23178 48473 5064 VDDPOST VDDPOST pch l=0.04u w=0.12u
m23179 5071 5066 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23180 VDDPOST 4935 5070 VDDPOST pch l=0.04u w=0.8u
m23181 5085 5094 48473 VDDPOST pch l=0.04u w=0.12u
m23182 5087 5248 5085 VDDPOST pch l=0.04u w=0.8u
m23183 5073 4671 5015 5014 pch l=0.04u w=0.4u
m23184 5074 4671 4 5014 pch l=0.04u w=0.4u
m23185 5075 4671 5015 5014 pch l=0.04u w=0.4u
m23186 5076 4671 4 5014 pch l=0.04u w=0.4u
m23187 5077 4671 5015 5014 pch l=0.04u w=0.4u
m23188 5078 4671 4 5014 pch l=0.04u w=0.4u
m23189 5079 4671 5015 5014 pch l=0.04u w=0.4u
m23190 5080 4671 4 5014 pch l=0.04u w=0.4u
m23191 5081 4671 5015 5014 pch l=0.04u w=0.4u
m23192 5082 4671 4 5014 pch l=0.04u w=0.4u
m23193 5083 4672 4 5014 pch l=0.04u w=0.4u
m23194 5084 4672 4 5014 pch l=0.04u w=0.4u
m23195 5088 5143 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23196 5089 4989 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23197 5090 5070 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23198 VSS 4573 5073 5014 pch l=0.04u w=0.4u
m23199 5015 4573 5074 5014 pch l=0.04u w=0.4u
m23200 VSS 4573 5075 5014 pch l=0.04u w=0.4u
m23201 5015 4573 5076 5014 pch l=0.04u w=0.4u
m23202 VSS 4573 5077 5014 pch l=0.04u w=0.4u
m23203 5015 4573 5078 5014 pch l=0.04u w=0.4u
m23204 VSS 4573 5079 5014 pch l=0.04u w=0.4u
m23205 5015 4573 5080 5014 pch l=0.04u w=0.4u
m23206 VSS 4573 5081 5014 pch l=0.04u w=0.4u
m23207 5015 4573 5082 5014 pch l=0.04u w=0.4u
m23208 5015 4574 5083 5014 pch l=0.04u w=0.4u
m23209 5015 4574 5084 5014 pch l=0.04u w=0.4u
m23210 VDDPOST 5065 5090 VDDPOST pch l=0.04u w=0.8u
m23211 5094 5248 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23212 FOUT2 5132 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23213 5096 4989 5071 VDDPOST pch l=0.04u w=0.8u
m23214 5090 5065 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23215 VDDPOST 5132 FOUT2 VDDPOST pch l=0.04u w=0.8u
m23216 48969 5089 5096 VDDPOST pch l=0.04u w=0.12u
m23217 VDDPOST 5070 5090 VDDPOST pch l=0.04u w=0.8u
m23218 FOUT2 5132 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23219 VDDPOST 5111 48969 VDDPOST pch l=0.04u w=0.12u
m23220 VDDPOST 5112 5087 VDDPOST pch l=0.04u w=0.8u
m23221 VDDPOST 5132 FOUT2 VDDPOST pch l=0.04u w=0.8u
m23222 5098 4432 5015 5014 pch l=0.04u w=0.4u
m23223 5099 4432 4 5014 pch l=0.04u w=0.4u
m23224 5100 4432 5015 5014 pch l=0.04u w=0.4u
m23225 5101 4432 4 5014 pch l=0.04u w=0.4u
m23226 5102 4432 5015 5014 pch l=0.04u w=0.4u
m23227 5103 4432 4 5014 pch l=0.04u w=0.4u
m23228 5104 4432 5015 5014 pch l=0.04u w=0.4u
m23229 5105 4432 4 5014 pch l=0.04u w=0.4u
m23230 5106 4432 5015 5014 pch l=0.04u w=0.4u
m23231 5107 4432 4 5014 pch l=0.04u w=0.4u
m23232 5108 4433 4 5014 pch l=0.04u w=0.4u
m23233 5109 4433 4 5014 pch l=0.04u w=0.4u
m23234 5111 5096 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23235 5113 4858 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23236 FOUT2 5132 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23237 VSS 4532 5098 5014 pch l=0.04u w=0.4u
m23238 5015 4532 5099 5014 pch l=0.04u w=0.4u
m23239 VSS 4532 5100 5014 pch l=0.04u w=0.4u
m23240 5015 4532 5101 5014 pch l=0.04u w=0.4u
m23241 VSS 4532 5102 5014 pch l=0.04u w=0.4u
m23242 5015 4532 5103 5014 pch l=0.04u w=0.4u
m23243 VSS 4532 5104 5014 pch l=0.04u w=0.4u
m23244 5015 4532 5105 5014 pch l=0.04u w=0.4u
m23245 VSS 4532 5106 5014 pch l=0.04u w=0.4u
m23246 5015 4532 5107 5014 pch l=0.04u w=0.4u
m23247 5015 4533 5108 5014 pch l=0.04u w=0.4u
m23248 5015 4533 5109 5014 pch l=0.04u w=0.4u
m23249 5112 5117 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23250 VDDPOST 5527 5113 VDDPOST pch l=0.04u w=0.8u
m23251 VDDPOST 5132 FOUT2 VDDPOST pch l=0.04u w=0.8u
m23252 5115 5089 5111 VDDPOST pch l=0.04u w=0.8u
m23253 VDDPOST 4999 5112 VDDPOST pch l=0.04u w=0.8u
m23254 5113 5527 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23255 FOUT2 5132 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23256 49357 4989 5115 VDDPOST pch l=0.04u w=0.12u
m23257 VDDPOST 5132 FOUT2 VDDPOST pch l=0.04u w=0.8u
m23258 VDDPOST 5133 49357 VDDPOST pch l=0.04u w=0.12u
m23259 VDDPOST 5135 5117 VDDPOST pch l=0.04u w=0.8u
m23260 5130 5113 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23261 5118 4671 5015 5014 pch l=0.04u w=0.4u
m23262 5119 4671 4 5014 pch l=0.04u w=0.4u
m23263 5120 4671 5015 5014 pch l=0.04u w=0.4u
m23264 5121 4671 4 5014 pch l=0.04u w=0.4u
m23265 5122 4671 5015 5014 pch l=0.04u w=0.4u
m23266 5123 4671 4 5014 pch l=0.04u w=0.4u
m23267 5124 4671 5015 5014 pch l=0.04u w=0.4u
m23268 5125 4671 4 5014 pch l=0.04u w=0.4u
m23269 5126 4671 5015 5014 pch l=0.04u w=0.4u
m23270 5127 4671 4 5014 pch l=0.04u w=0.4u
m23271 5128 4672 4 5014 pch l=0.04u w=0.4u
m23272 5129 4672 4 5014 pch l=0.04u w=0.4u
m23273 5133 5115 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23274 49522 5087 VDDPOST VDDPOST pch l=0.04u w=0.24u
m23275 VDDREF 5137 5116 VDDREF pch l=0.26u w=0.4u
m23276 VDDPOST 5162 5132 VDDPOST pch l=0.04u w=0.8u
m23277 VSS 4573 5118 5014 pch l=0.04u w=0.4u
m23278 5015 4573 5119 5014 pch l=0.04u w=0.4u
m23279 VSS 4573 5120 5014 pch l=0.04u w=0.4u
m23280 5015 4573 5121 5014 pch l=0.04u w=0.4u
m23281 VSS 4573 5122 5014 pch l=0.04u w=0.4u
m23282 5015 4573 5123 5014 pch l=0.04u w=0.4u
m23283 VSS 4573 5124 5014 pch l=0.04u w=0.4u
m23284 5015 4573 5125 5014 pch l=0.04u w=0.4u
m23285 VSS 4573 5126 5014 pch l=0.04u w=0.4u
m23286 5015 4573 5127 5014 pch l=0.04u w=0.4u
m23287 5015 4574 5128 5014 pch l=0.04u w=0.4u
m23288 5015 4574 5129 5014 pch l=0.04u w=0.4u
m23289 5135 5248 49522 VDDPOST pch l=0.04u w=0.24u
m23290 5136 5113 5090 VDDPOST pch l=0.04u w=0.8u
m23291 5132 5162 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23292 5138 5182 5135 VDDPOST pch l=0.04u w=0.8u
m23293 49692 5130 5136 VDDPOST pch l=0.04u w=0.12u
m23294 VDDREF 2427 5137 VDDREF pch l=0.04u w=0.8u
m23295 VDDPOST 4962 5132 VDDPOST pch l=0.04u w=0.8u
m23296 5140 4989 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23297 VDDPOST 5156 49692 VDDPOST pch l=0.04u w=0.12u
m23298 5142 5137 VDDREF VDDREF pch l=0.04u w=0.8u
m23299 5138 5163 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23300 5156 5136 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23301 VDDPOST 5160 5143 VDDPOST pch l=0.04u w=0.8u
m23302 5144 4510 5015 5014 pch l=0.04u w=0.4u
m23303 5145 4510 4 5014 pch l=0.04u w=0.4u
m23304 5146 4509 5015 5014 pch l=0.04u w=0.4u
m23305 5147 4509 4 5014 pch l=0.04u w=0.4u
m23306 5148 4432 5015 5014 pch l=0.04u w=0.4u
m23307 5149 4432 4 5014 pch l=0.04u w=0.4u
m23308 5150 4432 5015 5014 pch l=0.04u w=0.4u
m23309 5151 4432 4 5014 pch l=0.04u w=0.4u
m23310 5152 4432 5015 5014 pch l=0.04u w=0.4u
m23311 5153 4432 4 5014 pch l=0.04u w=0.4u
m23312 5154 4433 4 5014 pch l=0.04u w=0.4u
m23313 5155 4433 4 5014 pch l=0.04u w=0.4u
m23314 5157 4989 5133 VDDPOST pch l=0.04u w=0.8u
m23315 VDDPOST 4999 5138 VDDPOST pch l=0.04u w=0.8u
m23316 5160 5162 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23317 VSS 4558 5144 5014 pch l=0.04u w=0.4u
m23318 5015 4558 5145 5014 pch l=0.04u w=0.4u
m23319 VSS 4557 5146 5014 pch l=0.04u w=0.4u
m23320 5015 4557 5147 5014 pch l=0.04u w=0.4u
m23321 VSS 4532 5148 5014 pch l=0.04u w=0.4u
m23322 5015 4532 5149 5014 pch l=0.04u w=0.4u
m23323 VSS 4532 5150 5014 pch l=0.04u w=0.4u
m23324 5015 4532 5151 5014 pch l=0.04u w=0.4u
m23325 VSS 4532 5152 5014 pch l=0.04u w=0.4u
m23326 5015 4532 5153 5014 pch l=0.04u w=0.4u
m23327 5015 4533 5154 5014 pch l=0.04u w=0.4u
m23328 5015 4533 5155 5014 pch l=0.04u w=0.4u
m23329 49972 5140 5157 VDDPOST pch l=0.04u w=0.12u
m23330 49978 5138 VDDPOST VDDPOST pch l=0.04u w=0.12u
m23331 5161 5130 5156 VDDPOST pch l=0.04u w=0.8u
m23332 5159 5142 VDDREF VDDREF pch l=0.26u w=0.4u
m23333 VDDPOST 5164 49972 VDDPOST pch l=0.04u w=0.12u
m23334 5163 5182 49978 VDDPOST pch l=0.04u w=0.12u
m23335 50074 5113 5161 VDDPOST pch l=0.04u w=0.12u
m23336 5162 5204 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23337 5164 5157 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23338 4999 5248 5163 VDDPOST pch l=0.04u w=0.8u
m23339 VDDPOST 5177 50074 VDDPOST pch l=0.04u w=0.12u
m23340 VDDPOST 5180 5162 VDDPOST pch l=0.04u w=0.8u
m23341 5177 5161 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23342 5165 4698 5015 5014 pch l=0.04u w=0.4u
m23343 5166 4698 4 5014 pch l=0.04u w=0.4u
m23344 5167 4697 5015 5014 pch l=0.04u w=0.4u
m23345 5168 4697 4 5014 pch l=0.04u w=0.4u
m23346 5169 4671 5015 5014 pch l=0.04u w=0.4u
m23347 5170 4671 4 5014 pch l=0.04u w=0.4u
m23348 5171 4671 5015 5014 pch l=0.04u w=0.4u
m23349 5172 4671 4 5014 pch l=0.04u w=0.4u
m23350 5173 4671 5015 5014 pch l=0.04u w=0.4u
m23351 5174 4671 4 5014 pch l=0.04u w=0.4u
m23352 5175 4672 4 5014 pch l=0.04u w=0.4u
m23353 5176 4672 4 5014 pch l=0.04u w=0.4u
m23354 5181 5140 5164 VDDPOST pch l=0.04u w=0.8u
m23355 5182 5248 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23356 VDDPOST 5179 5180 VDDPOST pch l=0.04u w=0.8u
m23357 VSS 4648 5165 5014 pch l=0.04u w=0.4u
m23358 5015 4648 5166 5014 pch l=0.04u w=0.4u
m23359 VSS 4647 5167 5014 pch l=0.04u w=0.4u
m23360 5015 4647 5168 5014 pch l=0.04u w=0.4u
m23361 VSS 4573 5169 5014 pch l=0.04u w=0.4u
m23362 5015 4573 5170 5014 pch l=0.04u w=0.4u
m23363 VSS 4573 5171 5014 pch l=0.04u w=0.4u
m23364 5015 4573 5172 5014 pch l=0.04u w=0.4u
m23365 VSS 4573 5173 5014 pch l=0.04u w=0.4u
m23366 5015 4573 5174 5014 pch l=0.04u w=0.4u
m23367 5015 4574 5175 5014 pch l=0.04u w=0.4u
m23368 5015 4574 5176 5014 pch l=0.04u w=0.4u
m23369 50350 4989 5181 VDDPOST pch l=0.04u w=0.12u
m23370 VDDPOST 5189 50350 VDDPOST pch l=0.04u w=0.12u
m23371 5186 5186 VDDREF VDDREF pch l=0.04u w=1u
m23372 FOUT1PH180 5226 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23373 5188 5177 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23374 VDDPOST 5204 5184 VDDPOST pch l=0.04u w=0.8u
m23375 5189 5181 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23376 VDDPOST 5226 FOUT1PH180 VDDPOST pch l=0.04u w=0.8u
m23377 FOUT1PH180 5226 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23378 5203 4876 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23379 5191 4510 5015 5014 pch l=0.04u w=0.4u
m23380 5192 4510 4 5014 pch l=0.04u w=0.4u
m23381 5193 4509 5015 5014 pch l=0.04u w=0.4u
m23382 5194 4509 4 5014 pch l=0.04u w=0.4u
m23383 5195 4506 5015 5014 pch l=0.04u w=0.4u
m23384 5196 4506 4 5014 pch l=0.04u w=0.4u
m23385 5197 4432 5015 5014 pch l=0.04u w=0.4u
m23386 5198 4432 4 5014 pch l=0.04u w=0.4u
m23387 5199 4432 5015 5014 pch l=0.04u w=0.4u
m23388 5200 4432 4 5014 pch l=0.04u w=0.4u
m23389 5201 4433 4 5014 pch l=0.04u w=0.4u
m23390 5202 4433 4 5014 pch l=0.04u w=0.4u
m23391 VDDPOST 5226 FOUT1PH180 VDDPOST pch l=0.04u w=0.8u
m23392 VDDPOST 5188 5203 VDDPOST pch l=0.04u w=0.8u
m23393 VDDPOST 5210 5204 VDDPOST pch l=0.04u w=0.8u
m23394 VSS 4558 5191 5014 pch l=0.04u w=0.4u
m23395 5015 4558 5192 5014 pch l=0.04u w=0.4u
m23396 VSS 4557 5193 5014 pch l=0.04u w=0.4u
m23397 5015 4557 5194 5014 pch l=0.04u w=0.4u
m23398 VSS 4554 5195 5014 pch l=0.04u w=0.4u
m23399 5015 4554 5196 5014 pch l=0.04u w=0.4u
m23400 VSS 4532 5197 5014 pch l=0.04u w=0.4u
m23401 5015 4532 5198 5014 pch l=0.04u w=0.4u
m23402 VSS 4532 5199 5014 pch l=0.04u w=0.4u
m23403 5015 4532 5200 5014 pch l=0.04u w=0.4u
m23404 5015 4533 5201 5014 pch l=0.04u w=0.4u
m23405 5015 4533 5202 5014 pch l=0.04u w=0.4u
m23406 FOUT1PH180 5226 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23407 5203 5042 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23408 5207 4989 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23409 50820 5204 VDDPOST VDDPOST pch l=0.04u w=0.12u
m23410 VDDPOST 5226 FOUT1PH180 VDDPOST pch l=0.04u w=0.8u
m23411 50862 5230 5206 VDDREF pch l=0.04u w=0.44u
m23412 5210 5277 50820 VDDPOST pch l=0.04u w=0.12u
m23413 FOUT1PH180 5226 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23414 VDDREF 5206 5208 VDDREF pch l=0.04u w=0.8u
m23415 5212 POSTDIV2[0] VDDPOST VDDPOST pch l=0.04u w=0.12u
m23416 5211 4989 5189 VDDPOST pch l=0.04u w=0.8u
m23417 5213 5257 5210 VDDPOST pch l=0.04u w=0.8u
m23418 VDDREF 5185 50862 VDDREF pch l=0.2u w=0.44u
m23419 VDDPOST 5226 FOUT1PH180 VDDPOST pch l=0.04u w=0.8u
m23420 VDDPOST 5188 5212 VDDPOST pch l=0.04u w=0.4u
m23421 51067 5207 5211 VDDPOST pch l=0.04u w=0.12u
m23422 5214 4698 5015 5014 pch l=0.04u w=0.4u
m23423 5215 4698 4 5014 pch l=0.04u w=0.4u
m23424 5216 4697 5015 5014 pch l=0.04u w=0.4u
m23425 5217 4697 4 5014 pch l=0.04u w=0.4u
m23426 5218 4694 5015 5014 pch l=0.04u w=0.4u
m23427 5219 4694 4 5014 pch l=0.04u w=0.4u
m23428 5220 4671 5015 5014 pch l=0.04u w=0.4u
m23429 5221 4671 4 5014 pch l=0.04u w=0.4u
m23430 5222 4671 5015 5014 pch l=0.04u w=0.4u
m23431 5223 4671 4 5014 pch l=0.04u w=0.4u
m23432 5224 4672 4 5014 pch l=0.04u w=0.4u
m23433 5225 4672 4 5014 pch l=0.04u w=0.4u
m23434 5212 5188 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23435 5227 5230 VDDREF VDDREF pch l=0.04u w=0.8u
m23436 VDDPOST 5229 51067 VDDPOST pch l=0.04u w=0.12u
m23437 51135 5185 VDDREF VDDREF pch l=0.2u w=0.44u
m23438 VDDPOST 5233 5213 VDDPOST pch l=0.04u w=0.8u
m23439 VDDPOST 5343 5226 VDDPOST pch l=0.04u w=0.8u
m23440 VSS 4648 5214 5014 pch l=0.04u w=0.4u
m23441 5015 4648 5215 5014 pch l=0.04u w=0.4u
m23442 VSS 4647 5216 5014 pch l=0.04u w=0.4u
m23443 5015 4647 5217 5014 pch l=0.04u w=0.4u
m23444 VSS 4644 5218 5014 pch l=0.04u w=0.4u
m23445 5015 4644 5219 5014 pch l=0.04u w=0.4u
m23446 VSS 4573 5220 5014 pch l=0.04u w=0.4u
m23447 5015 4573 5221 5014 pch l=0.04u w=0.4u
m23448 VSS 4573 5222 5014 pch l=0.04u w=0.4u
m23449 5015 4573 5223 5014 pch l=0.04u w=0.4u
m23450 5015 4574 5224 5014 pch l=0.04u w=0.4u
m23451 5015 4574 5225 5014 pch l=0.04u w=0.4u
m23452 5229 5211 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23453 5230 5206 51135 VDDREF pch l=0.04u w=0.44u
m23454 51197 5213 VDDPOST VDDPOST pch l=0.04u w=0.12u
m23455 5226 5343 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23456 4935 5203 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23457 5233 5257 51197 VDDPOST pch l=0.04u w=0.12u
m23458 VDDPOST 5017 5226 VDDPOST pch l=0.04u w=0.8u
m23459 5235 5207 5229 VDDPOST pch l=0.04u w=0.8u
m23460 VDDPOST 5212 4935 VDDPOST pch l=0.04u w=0.8u
m23461 5232 5208 VDDREF VDDREF pch l=0.04u w=0.8u
m23462 5184 5277 5233 VDDPOST pch l=0.04u w=0.8u
m23463 51427 4989 5235 VDDPOST pch l=0.04u w=0.12u
m23464 4935 5439 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23465 VDDREF 5271 5232 VDDREF pch l=0.04u w=0.8u
m23466 VDDPOST 5253 5248 VDDPOST pch l=0.04u w=0.8u
m23467 5236 4510 5015 5014 pch l=0.04u w=0.4u
m23468 5237 4510 4 5014 pch l=0.04u w=0.4u
m23469 5238 4509 5015 5014 pch l=0.04u w=0.4u
m23470 5239 4509 4 5014 pch l=0.04u w=0.4u
m23471 5240 4508 5015 5014 pch l=0.04u w=0.4u
m23472 5241 4508 4 5014 pch l=0.04u w=0.4u
m23473 5242 4432 5015 5014 pch l=0.04u w=0.4u
m23474 5243 4432 4 5014 pch l=0.04u w=0.4u
m23475 5244 4432 5015 5014 pch l=0.04u w=0.4u
m23476 5245 4432 4 5014 pch l=0.04u w=0.4u
m23477 5246 4433 4 5014 pch l=0.04u w=0.4u
m23478 5247 4433 4 5014 pch l=0.04u w=0.4u
m23479 VDDPOST 5254 51427 VDDPOST pch l=0.04u w=0.12u
m23480 5253 5343 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23481 VSS 4558 5236 5014 pch l=0.04u w=0.4u
m23482 5015 4558 5237 5014 pch l=0.04u w=0.4u
m23483 VSS 4557 5238 5014 pch l=0.04u w=0.4u
m23484 5015 4557 5239 5014 pch l=0.04u w=0.4u
m23485 VSS 4556 5240 5014 pch l=0.04u w=0.4u
m23486 5015 4556 5241 5014 pch l=0.04u w=0.4u
m23487 VSS 4532 5242 5014 pch l=0.04u w=0.4u
m23488 5015 4532 5243 5014 pch l=0.04u w=0.4u
m23489 VSS 4532 5244 5014 pch l=0.04u w=0.4u
m23490 5015 4532 5245 5014 pch l=0.04u w=0.4u
m23491 5015 4533 5246 5014 pch l=0.04u w=0.4u
m23492 5015 4533 5247 5014 pch l=0.04u w=0.4u
m23493 5254 5235 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23494 4935 5203 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23495 5255 5277 5252 VDDPOST pch l=0.04u w=0.8u
m23496 51573 5274 5251 VDDREF pch l=0.04u w=0.44u
m23497 VDDPOST 5212 4935 VDDPOST pch l=0.04u w=0.8u
m23498 51632 5257 5255 VDDPOST pch l=0.04u w=0.12u
m23499 VDDREF 5251 5256 VDDREF pch l=0.04u w=0.8u
m23500 5257 5277 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23501 VDDREF 5185 51573 VDDREF pch l=0.2u w=0.44u
m23502 5038 5189 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23503 4935 5439 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23504 VDDPOST 5270 51632 VDDPOST pch l=0.04u w=0.12u
m23505 VDDPOST 5277 5257 VDDPOST pch l=0.04u w=0.8u
m23506 VDDPOST 5254 5038 VDDPOST pch l=0.04u w=0.8u
m23507 5270 5255 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23508 5271 5274 VDDREF VDDREF pch l=0.04u w=0.8u
m23509 51844 5185 VDDREF VDDREF pch l=0.2u w=0.44u
m23510 5257 5277 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23511 5258 4698 5015 5014 pch l=0.04u w=0.4u
m23512 5259 4698 4 5014 pch l=0.04u w=0.4u
m23513 5260 4697 5015 5014 pch l=0.04u w=0.4u
m23514 5261 4697 4 5014 pch l=0.04u w=0.4u
m23515 5262 4696 5015 5014 pch l=0.04u w=0.4u
m23516 5263 4696 4 5014 pch l=0.04u w=0.4u
m23517 5264 4671 5015 5014 pch l=0.04u w=0.4u
m23518 5265 4671 4 5014 pch l=0.04u w=0.4u
m23519 5266 4671 5015 5014 pch l=0.04u w=0.4u
m23520 5267 4671 4 5014 pch l=0.04u w=0.4u
m23521 5268 4672 4 5014 pch l=0.04u w=0.4u
m23522 5269 4672 4 5014 pch l=0.04u w=0.4u
m23523 5038 5254 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23524 5272 4858 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23525 5274 5251 51844 VDDREF pch l=0.04u w=0.44u
m23526 VDDPOST 5277 5257 VDDPOST pch l=0.04u w=0.8u
m23527 VSS 4648 5258 5014 pch l=0.04u w=0.4u
m23528 5015 4648 5259 5014 pch l=0.04u w=0.4u
m23529 VSS 4647 5260 5014 pch l=0.04u w=0.4u
m23530 5015 4647 5261 5014 pch l=0.04u w=0.4u
m23531 VSS 4646 5262 5014 pch l=0.04u w=0.4u
m23532 5015 4646 5263 5014 pch l=0.04u w=0.4u
m23533 VSS 4573 5264 5014 pch l=0.04u w=0.4u
m23534 5015 4573 5265 5014 pch l=0.04u w=0.4u
m23535 VSS 4573 5266 5014 pch l=0.04u w=0.4u
m23536 5015 4573 5267 5014 pch l=0.04u w=0.4u
m23537 5015 4574 5268 5014 pch l=0.04u w=0.4u
m23538 5015 4574 5269 5014 pch l=0.04u w=0.4u
m23539 VDDPOST 5189 5038 VDDPOST pch l=0.04u w=0.8u
m23540 5275 5257 5270 VDDPOST pch l=0.04u w=0.8u
m23541 52001 5277 5275 VDDPOST pch l=0.04u w=0.12u
m23542 5276 4858 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23543 5277 FOUT1PH180 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23544 5278 5229 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23545 VDDPOST 5291 52001 VDDPOST pch l=0.04u w=0.12u
m23546 VDDPOST 5177 5276 VDDPOST pch l=0.04u w=0.8u
m23547 VDDPOST FOUT1PH180 5277 VDDPOST pch l=0.04u w=0.8u
m23548 5291 5275 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23549 5277 FOUT1PH180 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23550 5279 4510 5015 5014 pch l=0.04u w=0.4u
m23551 5280 4510 4 5014 pch l=0.04u w=0.4u
m23552 5281 4509 5015 5014 pch l=0.04u w=0.4u
m23553 5282 4509 4 5014 pch l=0.04u w=0.4u
m23554 5283 4508 5015 5014 pch l=0.04u w=0.4u
m23555 5284 4508 4 5014 pch l=0.04u w=0.4u
m23556 5285 4432 5015 5014 pch l=0.04u w=0.4u
m23557 5286 4432 4 5014 pch l=0.04u w=0.4u
m23558 5287 4432 5015 5014 pch l=0.04u w=0.4u
m23559 5288 4432 4 5014 pch l=0.04u w=0.4u
m23560 5289 4433 4 5014 pch l=0.04u w=0.4u
m23561 5290 4433 4 5014 pch l=0.04u w=0.4u
m23562 5292 4977 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23563 5293 5272 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23564 VDDPOST FOUT1PH180 5277 VDDPOST pch l=0.04u w=0.8u
m23565 VSS 4558 5279 5014 pch l=0.04u w=0.4u
m23566 5015 4558 5280 5014 pch l=0.04u w=0.4u
m23567 VSS 4557 5281 5014 pch l=0.04u w=0.4u
m23568 5015 4557 5282 5014 pch l=0.04u w=0.4u
m23569 VSS 4556 5283 5014 pch l=0.04u w=0.4u
m23570 5015 4556 5284 5014 pch l=0.04u w=0.4u
m23571 VSS 4532 5285 5014 pch l=0.04u w=0.4u
m23572 5015 4532 5286 5014 pch l=0.04u w=0.4u
m23573 VSS 4532 5287 5014 pch l=0.04u w=0.4u
m23574 5015 4532 5288 5014 pch l=0.04u w=0.4u
m23575 5015 4533 5289 5014 pch l=0.04u w=0.4u
m23576 5015 4533 5290 5014 pch l=0.04u w=0.4u
m23577 VDDPOST 5278 5292 VDDPOST pch l=0.04u w=0.8u
m23578 5294 5291 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23579 VDDPOST 4935 5293 VDDPOST pch l=0.04u w=0.8u
m23580 5292 5254 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23581 5295 FOUTPOSTDIV VDDPOST VDDPOST pch l=0.04u w=0.8u
m23582 5252 5204 5291 VDDPOST pch l=0.04u w=0.8u
m23583 5297 5293 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23584 5310 4956 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23585 5204 5291 5252 VDDPOST pch l=0.04u w=0.8u
m23586 VDDPOST 5276 5297 VDDPOST pch l=0.04u w=0.8u
m23587 5311 5295 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23588 5298 4698 5015 5014 pch l=0.04u w=0.4u
m23589 5299 4698 4 5014 pch l=0.04u w=0.4u
m23590 5300 4697 5015 5014 pch l=0.04u w=0.4u
m23591 5301 4697 4 5014 pch l=0.04u w=0.4u
m23592 5302 4696 5015 5014 pch l=0.04u w=0.4u
m23593 5303 4696 4 5014 pch l=0.04u w=0.4u
m23594 5304 4671 5015 5014 pch l=0.04u w=0.4u
m23595 5305 4671 4 5014 pch l=0.04u w=0.4u
m23596 5306 4671 5015 5014 pch l=0.04u w=0.4u
m23597 5307 4671 4 5014 pch l=0.04u w=0.4u
m23598 5308 4672 4 5014 pch l=0.04u w=0.4u
m23599 5309 4672 4 5014 pch l=0.04u w=0.4u
m23600 VDDPOST 4708 5310 VDDPOST pch l=0.04u w=0.8u
m23601 5297 5276 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23602 VDDPOST 5295 5311 VDDPOST pch l=0.04u w=0.8u
m23603 VSS 4648 5298 5014 pch l=0.04u w=0.4u
m23604 5015 4648 5299 5014 pch l=0.04u w=0.4u
m23605 VSS 4647 5300 5014 pch l=0.04u w=0.4u
m23606 5015 4647 5301 5014 pch l=0.04u w=0.4u
m23607 VSS 4646 5302 5014 pch l=0.04u w=0.4u
m23608 5015 4646 5303 5014 pch l=0.04u w=0.4u
m23609 VSS 4573 5304 5014 pch l=0.04u w=0.4u
m23610 5015 4573 5305 5014 pch l=0.04u w=0.4u
m23611 VSS 4573 5306 5014 pch l=0.04u w=0.4u
m23612 5015 4573 5307 5014 pch l=0.04u w=0.4u
m23613 5015 4574 5308 5014 pch l=0.04u w=0.4u
m23614 5015 4574 5309 5014 pch l=0.04u w=0.4u
m23615 5310 4708 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23616 VDDPOST 5293 5297 VDDPOST pch l=0.04u w=0.8u
m23617 5318 5317 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23618 5320 5295 5319 VDDPOST pch l=0.04u w=0.8u
m23619 5321 5310 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23620 5322 5323 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23621 5324 5318 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23622 52943 5311 5320 VDDPOST pch l=0.04u w=0.12u
m23623 VDDPOST 5291 5324 VDDPOST pch l=0.04u w=0.8u
m23624 VDDPOST 5343 52943 VDDPOST pch l=0.04u w=0.12u
m23625 5325 4510 5015 5014 pch l=0.04u w=0.4u
m23626 5326 4510 4 5014 pch l=0.04u w=0.4u
m23627 5327 4509 5015 5014 pch l=0.04u w=0.4u
m23628 5328 4509 4 5014 pch l=0.04u w=0.4u
m23629 5329 4508 5015 5014 pch l=0.04u w=0.4u
m23630 5330 4508 4 5014 pch l=0.04u w=0.4u
m23631 5331 4432 5015 5014 pch l=0.04u w=0.4u
m23632 5332 4432 4 5014 pch l=0.04u w=0.4u
m23633 5333 4432 5015 5014 pch l=0.04u w=0.4u
m23634 5334 4432 4 5014 pch l=0.04u w=0.4u
m23635 5335 4433 4 5014 pch l=0.04u w=0.4u
m23636 5336 4433 4 5014 pch l=0.04u w=0.4u
m23637 5340 5310 5337 VDDPOST pch l=0.04u w=0.8u
m23638 5341 5322 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23639 5343 5320 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23640 VSS 4558 5325 5014 pch l=0.04u w=0.4u
m23641 5015 4558 5326 5014 pch l=0.04u w=0.4u
m23642 VSS 4557 5327 5014 pch l=0.04u w=0.4u
m23643 5015 4557 5328 5014 pch l=0.04u w=0.4u
m23644 VSS 4556 5329 5014 pch l=0.04u w=0.4u
m23645 5015 4556 5330 5014 pch l=0.04u w=0.4u
m23646 VSS 4532 5331 5014 pch l=0.04u w=0.4u
m23647 5015 4532 5332 5014 pch l=0.04u w=0.4u
m23648 VSS 4532 5333 5014 pch l=0.04u w=0.4u
m23649 5015 4532 5334 5014 pch l=0.04u w=0.4u
m23650 5015 4533 5335 5014 pch l=0.04u w=0.4u
m23651 5015 4533 5336 5014 pch l=0.04u w=0.4u
m23652 53128 5321 5340 VDDPOST pch l=0.04u w=0.12u
m23653 VDDPOST 5527 5341 VDDPOST pch l=0.04u w=0.8u
m23654 VDDPOST 5324 5342 VDDPOST pch l=0.04u w=0.8u
m23655 VDDPOST 5362 53128 VDDPOST pch l=0.04u w=0.12u
m23656 5341 5527 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23657 5361 5342 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23658 5362 5340 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23659 5363 5343 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23660 VDDPOST 5343 5363 VDDPOST pch l=0.04u w=0.8u
m23661 5377 5341 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23662 5378 5676 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23663 5365 4698 5015 5014 pch l=0.04u w=0.4u
m23664 5366 4698 4 5014 pch l=0.04u w=0.4u
m23665 5367 4697 5015 5014 pch l=0.04u w=0.4u
m23666 5368 4697 4 5014 pch l=0.04u w=0.4u
m23667 5369 4696 5015 5014 pch l=0.04u w=0.4u
m23668 5370 4696 4 5014 pch l=0.04u w=0.4u
m23669 5371 4671 5015 5014 pch l=0.04u w=0.4u
m23670 5372 4671 4 5014 pch l=0.04u w=0.4u
m23671 5373 4671 5015 5014 pch l=0.04u w=0.4u
m23672 5374 4671 4 5014 pch l=0.04u w=0.4u
m23673 5375 4672 4 5014 pch l=0.04u w=0.4u
m23674 5376 4672 4 5014 pch l=0.04u w=0.4u
m23675 5379 5321 5362 VDDPOST pch l=0.04u w=0.8u
m23676 VDDPOST 5324 5378 VDDPOST pch l=0.04u w=0.8u
m23677 VSS 4648 5365 5014 pch l=0.04u w=0.4u
m23678 5015 4648 5366 5014 pch l=0.04u w=0.4u
m23679 VSS 4647 5367 5014 pch l=0.04u w=0.4u
m23680 5015 4647 5368 5014 pch l=0.04u w=0.4u
m23681 VSS 4646 5369 5014 pch l=0.04u w=0.4u
m23682 5015 4646 5370 5014 pch l=0.04u w=0.4u
m23683 VSS 4573 5371 5014 pch l=0.04u w=0.4u
m23684 5015 4573 5372 5014 pch l=0.04u w=0.4u
m23685 VSS 4573 5373 5014 pch l=0.04u w=0.4u
m23686 5015 4573 5374 5014 pch l=0.04u w=0.4u
m23687 5015 4574 5375 5014 pch l=0.04u w=0.4u
m23688 5015 4574 5376 5014 pch l=0.04u w=0.4u
m23689 53512 5310 5379 VDDPOST pch l=0.04u w=0.12u
m23690 5392 5343 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23691 5378 5324 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23692 5393 5341 5297 VDDPOST pch l=0.04u w=0.8u
m23693 VDDPOST 5394 53512 VDDPOST pch l=0.04u w=0.12u
m23694 53601 5377 5393 VDDPOST pch l=0.04u w=0.12u
m23695 5394 5379 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23696 VDDPOST 5409 53601 VDDPOST pch l=0.04u w=0.12u
m23697 FOUT4 5378 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23698 5396 5311 5392 VDDPOST pch l=0.04u w=0.8u
m23699 5409 5393 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23700 VDDPOST 5378 FOUT4 VDDPOST pch l=0.04u w=0.8u
m23701 53816 5295 5396 VDDPOST pch l=0.04u w=0.12u
m23702 5397 4510 5015 5014 pch l=0.04u w=0.4u
m23703 5398 4510 4 5014 pch l=0.04u w=0.4u
m23704 5399 4509 5015 5014 pch l=0.04u w=0.4u
m23705 5400 4509 4 5014 pch l=0.04u w=0.4u
m23706 5401 4508 5015 5014 pch l=0.04u w=0.4u
m23707 5402 4508 4 5014 pch l=0.04u w=0.4u
m23708 5403 4432 5015 5014 pch l=0.04u w=0.4u
m23709 5404 4432 4 5014 pch l=0.04u w=0.4u
m23710 5405 4432 5015 5014 pch l=0.04u w=0.4u
m23711 5406 4432 4 5014 pch l=0.04u w=0.4u
m23712 5407 4433 4 5014 pch l=0.04u w=0.4u
m23713 5408 4433 4 5014 pch l=0.04u w=0.4u
m23714 FOUT4 5378 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23715 VDDPOST 5424 53816 VDDPOST pch l=0.04u w=0.12u
m23716 VSS 4558 5397 5014 pch l=0.04u w=0.4u
m23717 5015 4558 5398 5014 pch l=0.04u w=0.4u
m23718 VSS 4557 5399 5014 pch l=0.04u w=0.4u
m23719 5015 4557 5400 5014 pch l=0.04u w=0.4u
m23720 VSS 4556 5401 5014 pch l=0.04u w=0.4u
m23721 5015 4556 5402 5014 pch l=0.04u w=0.4u
m23722 VSS 4532 5403 5014 pch l=0.04u w=0.4u
m23723 5015 4532 5404 5014 pch l=0.04u w=0.4u
m23724 VSS 4532 5405 5014 pch l=0.04u w=0.4u
m23725 5015 4532 5406 5014 pch l=0.04u w=0.4u
m23726 5015 4533 5407 5014 pch l=0.04u w=0.4u
m23727 5015 4533 5408 5014 pch l=0.04u w=0.4u
m23728 5410 5310 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23729 VDDPOST 5378 FOUT4 VDDPOST pch l=0.04u w=0.8u
m23730 5423 5377 5409 VDDPOST pch l=0.04u w=0.8u
m23731 5424 5396 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23732 FOUT4 5378 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23733 54064 5341 5423 VDDPOST pch l=0.04u w=0.12u
m23734 5425 5310 5394 VDDPOST pch l=0.04u w=0.8u
m23735 VDDPOST 5378 FOUT4 VDDPOST pch l=0.04u w=0.8u
m23736 VDDPOST 5439 54064 VDDPOST pch l=0.04u w=0.12u
m23737 5426 5424 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23738 54261 5410 5425 VDDPOST pch l=0.04u w=0.12u
m23739 FOUT4 5378 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23740 5439 5423 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23741 VDDPOST 5424 5426 VDDPOST pch l=0.04u w=0.8u
m23742 VDDPOST 5440 54261 VDDPOST pch l=0.04u w=0.12u
m23743 VDDPOST 5378 FOUT4 VDDPOST pch l=0.04u w=0.8u
m23744 5427 4698 5015 5014 pch l=0.04u w=0.4u
m23745 5428 4698 4 5014 pch l=0.04u w=0.4u
m23746 5429 4697 5015 5014 pch l=0.04u w=0.4u
m23747 5430 4697 4 5014 pch l=0.04u w=0.4u
m23748 5431 4696 5015 5014 pch l=0.04u w=0.4u
m23749 5432 4696 4 5014 pch l=0.04u w=0.4u
m23750 5433 4671 5015 5014 pch l=0.04u w=0.4u
m23751 5434 4671 4 5014 pch l=0.04u w=0.4u
m23752 5435 4671 5015 5014 pch l=0.04u w=0.4u
m23753 5436 4671 4 5014 pch l=0.04u w=0.4u
m23754 5437 4672 4 5014 pch l=0.04u w=0.4u
m23755 5438 4672 4 5014 pch l=0.04u w=0.4u
m23756 5440 5425 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23757 VSS 4648 5427 5014 pch l=0.04u w=0.4u
m23758 5015 4648 5428 5014 pch l=0.04u w=0.4u
m23759 VSS 4647 5429 5014 pch l=0.04u w=0.4u
m23760 5015 4647 5430 5014 pch l=0.04u w=0.4u
m23761 VSS 4646 5431 5014 pch l=0.04u w=0.4u
m23762 5015 4646 5432 5014 pch l=0.04u w=0.4u
m23763 VSS 4573 5433 5014 pch l=0.04u w=0.4u
m23764 5015 4573 5434 5014 pch l=0.04u w=0.4u
m23765 VSS 4573 5435 5014 pch l=0.04u w=0.4u
m23766 5015 4573 5436 5014 pch l=0.04u w=0.4u
m23767 5015 4574 5437 5014 pch l=0.04u w=0.4u
m23768 5015 4574 5438 5014 pch l=0.04u w=0.4u
m23769 5455 5424 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23770 5456 POSTDIV2[0] VDDPOST VDDPOST pch l=0.04u w=0.12u
m23771 VDDPOST 5361 5454 VDDPOST pch l=0.04u w=0.8u
m23772 VDDPOST 5409 5456 VDDPOST pch l=0.04u w=0.4u
m23773 5457 5410 5440 VDDPOST pch l=0.04u w=0.8u
m23774 5319 5455 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23775 5456 5409 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23776 54963 5310 5457 VDDPOST pch l=0.04u w=0.12u
m23777 5471 5361 5458 VDDPOST pch l=0.04u w=0.8u
m23778 VDDPOST 5473 54963 VDDPOST pch l=0.04u w=0.12u
m23779 5459 4510 5015 5014 pch l=0.04u w=0.4u
m23780 5460 4510 4 5014 pch l=0.04u w=0.4u
m23781 5461 4509 5015 5014 pch l=0.04u w=0.4u
m23782 5462 4509 4 5014 pch l=0.04u w=0.4u
m23783 5463 4507 5015 5014 pch l=0.04u w=0.4u
m23784 5464 4507 4 5014 pch l=0.04u w=0.4u
m23785 5465 4432 5015 5014 pch l=0.04u w=0.4u
m23786 5466 4432 4 5014 pch l=0.04u w=0.4u
m23787 5467 4432 5015 5014 pch l=0.04u w=0.4u
m23788 5468 4432 4 5014 pch l=0.04u w=0.4u
m23789 5469 4433 4 5014 pch l=0.04u w=0.4u
m23790 5470 4433 4 5014 pch l=0.04u w=0.4u
m23791 55218 5454 5471 VDDPOST pch l=0.04u w=0.12u
m23792 5472 FOUT1PH90 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23793 5473 5457 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23794 VSS 4558 5459 5014 pch l=0.04u w=0.4u
m23795 5015 4558 5460 5014 pch l=0.04u w=0.4u
m23796 VSS 4557 5461 5014 pch l=0.04u w=0.4u
m23797 5015 4557 5462 5014 pch l=0.04u w=0.4u
m23798 VSS 4555 5463 5014 pch l=0.04u w=0.4u
m23799 5015 4555 5464 5014 pch l=0.04u w=0.4u
m23800 VSS 4532 5465 5014 pch l=0.04u w=0.4u
m23801 5015 4532 5466 5014 pch l=0.04u w=0.4u
m23802 VSS 4532 5467 5014 pch l=0.04u w=0.4u
m23803 5015 4532 5468 5014 pch l=0.04u w=0.4u
m23804 5015 4533 5469 5014 pch l=0.04u w=0.4u
m23805 5015 4533 5470 5014 pch l=0.04u w=0.4u
m23806 VDDPOST 5487 55218 VDDPOST pch l=0.04u w=0.12u
m23807 5486 5456 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23808 VDDPOST FOUT1PH90 5472 VDDPOST pch l=0.04u w=0.8u
m23809 5487 5458 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23810 VDDPOST 5439 5486 VDDPOST pch l=0.04u w=0.8u
m23811 5472 FOUT1PH90 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23812 VDDPOST 5471 5487 VDDPOST pch l=0.04u w=0.8u
m23813 VDDPOST FOUT1PH90 5472 VDDPOST pch l=0.04u w=0.8u
m23814 5503 5310 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23815 5504 5486 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23816 5508 5454 5487 VDDPOST pch l=0.04u w=0.8u
m23817 5491 4698 5015 5014 pch l=0.04u w=0.4u
m23818 5492 4698 4 5014 pch l=0.04u w=0.4u
m23819 5493 4697 5015 5014 pch l=0.04u w=0.4u
m23820 5494 4697 4 5014 pch l=0.04u w=0.4u
m23821 5495 4695 5015 5014 pch l=0.04u w=0.4u
m23822 5496 4695 4 5014 pch l=0.04u w=0.4u
m23823 5497 4671 5015 5014 pch l=0.04u w=0.4u
m23824 5498 4671 4 5014 pch l=0.04u w=0.4u
m23825 5499 4671 5015 5014 pch l=0.04u w=0.4u
m23826 5500 4671 4 5014 pch l=0.04u w=0.4u
m23827 5501 4672 4 5014 pch l=0.04u w=0.4u
m23828 5502 4672 4 5014 pch l=0.04u w=0.4u
m23829 VDDPOST 5486 5504 VDDPOST pch l=0.04u w=0.8u
m23830 VDDPOST 5426 5505 VDDPOST pch l=0.04u w=0.8u
m23831 56093 5361 5508 VDDPOST pch l=0.04u w=0.24u
m23832 VSS 4648 5491 5014 pch l=0.04u w=0.4u
m23833 5015 4648 5492 5014 pch l=0.04u w=0.4u
m23834 VSS 4647 5493 5014 pch l=0.04u w=0.4u
m23835 5015 4647 5494 5014 pch l=0.04u w=0.4u
m23836 VSS 4645 5495 5014 pch l=0.04u w=0.4u
m23837 5015 4645 5496 5014 pch l=0.04u w=0.4u
m23838 VSS 4573 5497 5014 pch l=0.04u w=0.4u
m23839 5015 4573 5498 5014 pch l=0.04u w=0.4u
m23840 VSS 4573 5499 5014 pch l=0.04u w=0.4u
m23841 5015 4573 5500 5014 pch l=0.04u w=0.4u
m23842 5015 4574 5501 5014 pch l=0.04u w=0.4u
m23843 5015 4574 5502 5014 pch l=0.04u w=0.4u
m23844 5512 5310 5473 VDDPOST pch l=0.04u w=0.8u
m23845 5525 5505 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23846 VDDPOST 5564 56093 VDDPOST pch l=0.04u w=0.24u
m23847 56198 5503 5512 VDDPOST pch l=0.04u w=0.12u
m23848 5527 5549 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23849 5528 5792 5526 VDDREF pch l=0.1u w=1u
m23850 5531 5508 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23851 VDDPOST 5534 56198 VDDPOST pch l=0.04u w=0.12u
m23852 VDDPOST 5549 5527 VDDPOST pch l=0.04u w=0.8u
m23853 5533 5794 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23854 5526 5792 5528 VDDREF pch l=0.1u w=1u
m23855 5534 5512 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23856 VDDPOST 5426 5533 VDDPOST pch l=0.04u w=0.8u
m23857 5548 5458 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23858 5535 4510 5015 5014 pch l=0.04u w=0.4u
m23859 5536 4510 4 5014 pch l=0.04u w=0.4u
m23860 5537 4509 5015 5014 pch l=0.04u w=0.4u
m23861 5538 4509 4 5014 pch l=0.04u w=0.4u
m23862 5539 4507 5015 5014 pch l=0.04u w=0.4u
m23863 5540 4507 4 5014 pch l=0.04u w=0.4u
m23864 5541 4432 5015 5014 pch l=0.04u w=0.4u
m23865 5542 4432 4 5014 pch l=0.04u w=0.4u
m23866 5543 4432 5015 5014 pch l=0.04u w=0.4u
m23867 5544 4432 4 5014 pch l=0.04u w=0.4u
m23868 5545 4433 4 5014 pch l=0.04u w=0.4u
m23869 5546 4433 4 5014 pch l=0.04u w=0.4u
m23870 5549 4710 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23871 5533 5426 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23872 VDDPOST 5531 5548 VDDPOST pch l=0.04u w=0.8u
m23873 5550 5503 5534 VDDPOST pch l=0.04u w=0.8u
m23874 VSS 4558 5535 5014 pch l=0.04u w=0.4u
m23875 5015 4558 5536 5014 pch l=0.04u w=0.4u
m23876 VSS 4557 5537 5014 pch l=0.04u w=0.4u
m23877 5015 4557 5538 5014 pch l=0.04u w=0.4u
m23878 VSS 4555 5539 5014 pch l=0.04u w=0.4u
m23879 5015 4555 5540 5014 pch l=0.04u w=0.4u
m23880 VSS 4532 5541 5014 pch l=0.04u w=0.4u
m23881 5015 4532 5542 5014 pch l=0.04u w=0.4u
m23882 VSS 4532 5543 5014 pch l=0.04u w=0.4u
m23883 5015 4532 5544 5014 pch l=0.04u w=0.4u
m23884 5015 4533 5545 5014 pch l=0.04u w=0.4u
m23885 5015 4533 5546 5014 pch l=0.04u w=0.4u
m23886 VDDPOST 5767 5549 VDDPOST pch l=0.04u w=0.8u
m23887 56573 5783 VDDREF VDDREF pch l=0.25u w=1u
m23888 56604 5310 5550 VDDPOST pch l=0.04u w=0.12u
m23889 5549 5580 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23890 FOUT1PH90 5533 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23891 VDDPOST 5566 56604 VDDPOST pch l=0.04u w=0.12u
m23892 5564 5548 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23893 VDDPOST 5533 FOUT1PH90 VDDPOST pch l=0.04u w=0.8u
m23894 5526 5783 56573 VDDREF pch l=0.25u w=1u
m23895 5566 5550 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23896 5580 4715 VDDPOST VDDPOST pch l=0.04u w=0.12u
m23897 FOUT1PH90 5533 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23898 5567 4698 5015 5014 pch l=0.04u w=0.4u
m23899 5568 4698 4 5014 pch l=0.04u w=0.4u
m23900 5569 4697 5015 5014 pch l=0.04u w=0.4u
m23901 5570 4697 4 5014 pch l=0.04u w=0.4u
m23902 5571 4695 5015 5014 pch l=0.04u w=0.4u
m23903 5572 4695 4 5014 pch l=0.04u w=0.4u
m23904 5573 4671 5015 5014 pch l=0.04u w=0.4u
m23905 5574 4671 4 5014 pch l=0.04u w=0.4u
m23906 5575 4671 5015 5014 pch l=0.04u w=0.4u
m23907 5576 4671 4 5014 pch l=0.04u w=0.4u
m23908 5577 4672 4 5014 pch l=0.04u w=0.4u
m23909 5578 4672 4 5014 pch l=0.04u w=0.4u
m23910 VDDPOST 4708 5580 VDDPOST pch l=0.04u w=0.4u
m23911 VDDPOST 5361 5579 VDDPOST pch l=0.04u w=0.8u
m23912 56891 5783 5526 VDDREF pch l=0.25u w=1u
m23913 VDDPOST 5533 FOUT1PH90 VDDPOST pch l=0.04u w=0.8u
m23914 5594 POSTDIV1[0] VDDPOST VDDPOST pch l=0.04u w=0.12u
m23915 VSS 4648 5567 5014 pch l=0.04u w=0.4u
m23916 5015 4648 5568 5014 pch l=0.04u w=0.4u
m23917 VSS 4647 5569 5014 pch l=0.04u w=0.4u
m23918 5015 4647 5570 5014 pch l=0.04u w=0.4u
m23919 VSS 4645 5571 5014 pch l=0.04u w=0.4u
m23920 5015 4645 5572 5014 pch l=0.04u w=0.4u
m23921 VSS 4573 5573 5014 pch l=0.04u w=0.4u
m23922 5015 4573 5574 5014 pch l=0.04u w=0.4u
m23923 VSS 4573 5575 5014 pch l=0.04u w=0.4u
m23924 5015 4573 5576 5014 pch l=0.04u w=0.4u
m23925 5015 4574 5577 5014 pch l=0.04u w=0.4u
m23926 5015 4574 5578 5014 pch l=0.04u w=0.4u
m23927 5580 4708 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23928 FOUT1PH90 5533 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23929 VDDPOST 5534 5594 VDDPOST pch l=0.04u w=0.4u
m23930 VDDREF 5783 56891 VDDREF pch l=0.25u w=1u
m23931 5596 5361 5564 VDDPOST pch l=0.04u w=0.8u
m23932 VDDPOST 5533 FOUT1PH90 VDDPOST pch l=0.04u w=0.8u
m23933 5594 5534 VDDPOST VDDPOST pch l=0.04u w=0.4u
m23934 57115 5579 5596 VDDPOST pch l=0.04u w=0.12u
m23935 FOUT1PH90 5533 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23936 5597 4860 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23937 57171 5783 VDDREF VDDREF pch l=0.25u w=1u
m23938 VDDPOST 5612 57115 VDDPOST pch l=0.04u w=0.12u
m23939 VDDPOST 5533 FOUT1PH90 VDDPOST pch l=0.04u w=0.8u
m23940 5598 4433 4 5014 pch l=0.04u w=0.4u
m23941 5599 4433 4 5014 pch l=0.04u w=0.4u
m23942 5600 4433 4 5014 pch l=0.04u w=0.4u
m23943 5601 4433 4 5014 pch l=0.04u w=0.4u
m23944 5602 4433 4 5014 pch l=0.04u w=0.4u
m23945 5603 4433 4 5014 pch l=0.04u w=0.4u
m23946 5604 4433 4 5014 pch l=0.04u w=0.4u
m23947 5605 4433 4 5014 pch l=0.04u w=0.4u
m23948 5606 4433 4 5014 pch l=0.04u w=0.4u
m23949 5607 4433 4 5014 pch l=0.04u w=0.4u
m23950 5608 4433 4 5014 pch l=0.04u w=0.4u
m23951 5609 4433 4 5014 pch l=0.04u w=0.4u
m23952 5611 4956 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23953 5612 5458 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23954 5614 4860 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23955 5526 5783 57171 VDDREF pch l=0.25u w=1u
m23956 5015 4533 5598 5014 pch l=0.04u w=0.4u
m23957 5015 4533 5599 5014 pch l=0.04u w=0.4u
m23958 5015 4533 5600 5014 pch l=0.04u w=0.4u
m23959 5015 4533 5601 5014 pch l=0.04u w=0.4u
m23960 5015 4533 5602 5014 pch l=0.04u w=0.4u
m23961 5015 4533 5603 5014 pch l=0.04u w=0.4u
m23962 5015 4533 5604 5014 pch l=0.04u w=0.4u
m23963 5015 4533 5605 5014 pch l=0.04u w=0.4u
m23964 5015 4533 5606 5014 pch l=0.04u w=0.4u
m23965 5015 4533 5607 5014 pch l=0.04u w=0.4u
m23966 5015 4533 5608 5014 pch l=0.04u w=0.4u
m23967 5015 4533 5609 5014 pch l=0.04u w=0.4u
m23968 VDDPOST 5594 5611 VDDPOST pch l=0.04u w=0.8u
m23969 VDDPOST 5596 5612 VDDPOST pch l=0.04u w=0.8u
m23970 VDDPOST 5525 5613 VDDPOST pch l=0.04u w=0.8u
m23971 VDDPOST 4707 5614 VDDPOST pch l=0.04u w=0.8u
m23972 5611 5566 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23973 57451 5783 5526 VDDREF pch l=0.25u w=1u
m23974 5628 5579 5612 VDDPOST pch l=0.04u w=0.8u
m23975 5629 5525 5627 VDDPOST pch l=0.04u w=0.8u
m23976 5630 5597 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23977 VDDPOST 5566 5337 VDDPOST pch l=0.04u w=0.8u
m23978 57606 5361 5628 VDDPOST pch l=0.04u w=0.24u
m23979 VDDREF 5783 57451 VDDREF pch l=0.25u w=1u
m23980 57621 5613 5629 VDDPOST pch l=0.04u w=0.12u
m23981 VDDPOST 5504 5630 VDDPOST pch l=0.04u w=0.8u
m23982 5631 4672 4 5014 pch l=0.04u w=0.4u
m23983 5632 4672 4 5014 pch l=0.04u w=0.4u
m23984 5633 4672 4 5014 pch l=0.04u w=0.4u
m23985 5634 4672 4 5014 pch l=0.04u w=0.4u
m23986 5635 4672 4 5014 pch l=0.04u w=0.4u
m23987 5636 4672 4 5014 pch l=0.04u w=0.4u
m23988 5637 4672 4 5014 pch l=0.04u w=0.4u
m23989 5638 4672 4 5014 pch l=0.04u w=0.4u
m23990 5639 4672 4 5014 pch l=0.04u w=0.4u
m23991 5640 4672 4 5014 pch l=0.04u w=0.4u
m23992 5641 4672 4 5014 pch l=0.04u w=0.4u
m23993 5642 4672 4 5014 pch l=0.04u w=0.4u
m23994 5337 5660 VDDPOST VDDPOST pch l=0.04u w=0.8u
m23995 VDDPOST 5676 57606 VDDPOST pch l=0.04u w=0.24u
m23996 VDDPOST 5657 57621 VDDPOST pch l=0.04u w=0.12u
m23997 57761 5783 VDDREF VDDREF pch l=0.25u w=1u
m23998 5015 4574 5631 5014 pch l=0.04u w=0.4u
m23999 5015 4574 5632 5014 pch l=0.04u w=0.4u
m24000 5015 4574 5633 5014 pch l=0.04u w=0.4u
m24001 5015 4574 5634 5014 pch l=0.04u w=0.4u
m24002 5015 4574 5635 5014 pch l=0.04u w=0.4u
m24003 5015 4574 5636 5014 pch l=0.04u w=0.4u
m24004 5015 4574 5637 5014 pch l=0.04u w=0.4u
m24005 5015 4574 5638 5014 pch l=0.04u w=0.4u
m24006 5015 4574 5639 5014 pch l=0.04u w=0.4u
m24007 5015 4574 5640 5014 pch l=0.04u w=0.4u
m24008 5015 4574 5641 5014 pch l=0.04u w=0.4u
m24009 5015 4574 5642 5014 pch l=0.04u w=0.4u
m24010 VDDPOST 5693 5337 VDDPOST pch l=0.04u w=0.8u
m24011 5644 5628 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24012 5657 5627 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24013 5658 5630 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24014 VDDPOST 5629 5657 VDDPOST pch l=0.04u w=0.8u
m24015 VDDPOST 5614 5658 VDDPOST pch l=0.04u w=0.8u
m24016 5511 5783 57761 VDDREF pch l=0.25u w=1u
m24017 5661 5458 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24018 VDDPOST 5690 5660 VDDPOST pch l=0.04u w=0.4u
m24019 5658 5614 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24020 VDDPOST 5644 5661 VDDPOST pch l=0.04u w=0.8u
m24021 5675 5613 5657 VDDPOST pch l=0.04u w=0.8u
m24022 5660 5690 VDDPOST VDDPOST pch l=0.04u w=0.4u
m24023 VDDPOST 5630 5658 VDDPOST pch l=0.04u w=0.8u
m24024 58087 5783 5511 VDDREF pch l=0.25u w=1u
m24025 5663 4433 4 5014 pch l=0.04u w=0.4u
m24026 5664 4433 4 5014 pch l=0.04u w=0.4u
m24027 5665 4433 4 5014 pch l=0.04u w=0.4u
m24028 5666 4433 4 5014 pch l=0.04u w=0.4u
m24029 5667 4433 4 5014 pch l=0.04u w=0.4u
m24030 5668 4433 4 5014 pch l=0.04u w=0.4u
m24031 5669 4433 4 5014 pch l=0.04u w=0.4u
m24032 5670 4433 4 5014 pch l=0.04u w=0.4u
m24033 5671 4433 4 5014 pch l=0.04u w=0.4u
m24034 5672 4433 4 5014 pch l=0.04u w=0.4u
m24035 5673 4433 4 5014 pch l=0.04u w=0.4u
m24036 5674 4433 4 5014 pch l=0.04u w=0.4u
m24037 58115 5525 5675 VDDPOST pch l=0.04u w=0.24u
m24038 VDDPOST POSTDIV1[0] 5660 VDDPOST pch l=0.04u w=0.12u
m24039 5015 4533 5663 5014 pch l=0.04u w=0.4u
m24040 5015 4533 5664 5014 pch l=0.04u w=0.4u
m24041 5015 4533 5665 5014 pch l=0.04u w=0.4u
m24042 5015 4533 5666 5014 pch l=0.04u w=0.4u
m24043 5015 4533 5667 5014 pch l=0.04u w=0.4u
m24044 5015 4533 5668 5014 pch l=0.04u w=0.4u
m24045 5015 4533 5669 5014 pch l=0.04u w=0.4u
m24046 5015 4533 5670 5014 pch l=0.04u w=0.4u
m24047 5015 4533 5671 5014 pch l=0.04u w=0.4u
m24048 5015 4533 5672 5014 pch l=0.04u w=0.4u
m24049 5015 4533 5673 5014 pch l=0.04u w=0.4u
m24050 5015 4533 5674 5014 pch l=0.04u w=0.4u
m24051 5676 5661 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24052 VDDPOST 5724 58115 VDDPOST pch l=0.04u w=0.24u
m24053 VDDREF 5783 58087 VDDREF pch l=0.25u w=1u
m24054 5689 4711 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24055 5691 5675 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24056 VDDPOST 5473 5690 VDDPOST pch l=0.04u w=0.8u
m24057 58381 5783 VDDREF VDDREF pch l=0.25u w=1u
m24058 5692 4711 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24059 5706 5627 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24060 VDDPOST 4953 5458 VDDPOST pch l=0.04u w=0.8u
m24061 VDDPOST 5767 5692 VDDPOST pch l=0.04u w=0.8u
m24062 VDDPOST 5394 5693 VDDPOST pch l=0.04u w=0.8u
m24063 5511 5783 58381 VDDREF pch l=0.25u w=1u
m24064 VDDPOST 5691 5706 VDDPOST pch l=0.04u w=0.8u
m24065 5694 4672 4 5014 pch l=0.04u w=0.4u
m24066 5695 4672 4 5014 pch l=0.04u w=0.4u
m24067 5696 4672 4 5014 pch l=0.04u w=0.4u
m24068 5697 4672 4 5014 pch l=0.04u w=0.4u
m24069 5698 4672 4 5014 pch l=0.04u w=0.4u
m24070 5699 4672 4 5014 pch l=0.04u w=0.4u
m24071 5700 4672 4 5014 pch l=0.04u w=0.4u
m24072 5701 4672 4 5014 pch l=0.04u w=0.4u
m24073 5702 4672 4 5014 pch l=0.04u w=0.4u
m24074 5703 4672 4 5014 pch l=0.04u w=0.4u
m24075 5704 4672 4 5014 pch l=0.04u w=0.4u
m24076 5705 4672 4 5014 pch l=0.04u w=0.4u
m24077 5693 5690 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24078 5015 4574 5694 5014 pch l=0.04u w=0.4u
m24079 5015 4574 5695 5014 pch l=0.04u w=0.4u
m24080 5015 4574 5696 5014 pch l=0.04u w=0.4u
m24081 5015 4574 5697 5014 pch l=0.04u w=0.4u
m24082 5015 4574 5698 5014 pch l=0.04u w=0.4u
m24083 5015 4574 5699 5014 pch l=0.04u w=0.4u
m24084 5015 4574 5700 5014 pch l=0.04u w=0.4u
m24085 5015 4574 5701 5014 pch l=0.04u w=0.4u
m24086 5015 4574 5702 5014 pch l=0.04u w=0.4u
m24087 5015 4574 5703 5014 pch l=0.04u w=0.4u
m24088 5015 4574 5704 5014 pch l=0.04u w=0.4u
m24089 5015 4574 5705 5014 pch l=0.04u w=0.4u
m24090 VDDPOST 4965 5693 VDDPOST pch l=0.04u w=0.8u
m24091 5721 5689 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24092 5722 5257 5708 VDDPOST pch l=0.04u w=0.8u
m24093 58662 5783 5511 VDDREF pch l=0.25u w=1u
m24094 5724 5706 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24095 VDDPOST 5658 5721 VDDPOST pch l=0.04u w=0.8u
m24096 58702 5277 5722 VDDPOST pch l=0.04u w=0.12u
m24097 5727 5292 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24098 VDDPOST 5731 58702 VDDPOST pch l=0.04u w=0.12u
m24099 VDDREF 5783 58662 VDDREF pch l=0.25u w=1u
m24100 VDDPOST 5611 5727 VDDPOST pch l=0.04u w=0.8u
m24101 5730 5721 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24102 5731 5722 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24103 VDDPOST 5525 5728 VDDPOST pch l=0.04u w=0.8u
m24104 5014 4389 4 5014 pch l=0.04u w=0.4u
m24105 5014 4389 4 5014 pch l=0.04u w=0.4u
m24106 5014 4389 4 5014 pch l=0.04u w=0.4u
m24107 5014 4389 4 5014 pch l=0.04u w=0.4u
m24108 5014 4389 4 5014 pch l=0.04u w=0.4u
m24109 5014 4389 4 5014 pch l=0.04u w=0.4u
m24110 5014 4389 4 5014 pch l=0.04u w=0.4u
m24111 5014 4389 4 5014 pch l=0.04u w=0.4u
m24112 5014 4389 4 5014 pch l=0.04u w=0.4u
m24113 5014 4389 4 5014 pch l=0.04u w=0.4u
m24114 5014 4389 4 5014 pch l=0.04u w=0.4u
m24115 5014 4389 4 5014 pch l=0.04u w=0.4u
m24116 5727 5798 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24117 VDDPOST 5692 5730 VDDPOST pch l=0.04u w=0.8u
m24118 5732 5792 5511 VDDREF pch l=0.1u w=1u
m24119 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24120 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24121 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24122 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24123 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24124 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24125 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24126 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24127 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24128 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24129 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24130 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24131 5730 5692 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24132 5746 5277 5731 VDDPOST pch l=0.04u w=0.8u
m24133 5747 5525 5724 VDDPOST pch l=0.04u w=0.8u
m24134 5511 5792 5732 VDDREF pch l=0.1u w=1u
m24135 VDDPOST 5721 5730 VDDPOST pch l=0.04u w=0.8u
m24136 5748 5727 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24137 59106 5257 5746 VDDPOST pch l=0.04u w=0.12u
m24138 59107 5728 5747 VDDPOST pch l=0.04u w=0.12u
m24139 VDDPOST 5750 59106 VDDPOST pch l=0.04u w=0.12u
m24140 VDDPOST 5751 59107 VDDPOST pch l=0.04u w=0.12u
m24141 5749 4791 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24142 5750 5746 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24143 5751 5627 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24144 5752 5748 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24145 5014 4389 4 5014 pch l=0.04u w=0.4u
m24146 5014 4389 4 5014 pch l=0.04u w=0.4u
m24147 5014 4389 4 5014 pch l=0.04u w=0.4u
m24148 5014 4389 4 5014 pch l=0.04u w=0.4u
m24149 5014 4389 4 5014 pch l=0.04u w=0.4u
m24150 5014 4389 4 5014 pch l=0.04u w=0.4u
m24151 5014 4389 4 5014 pch l=0.04u w=0.4u
m24152 5014 4389 4 5014 pch l=0.04u w=0.4u
m24153 5014 4389 4 5014 pch l=0.04u w=0.4u
m24154 5014 4389 4 5014 pch l=0.04u w=0.4u
m24155 5014 4389 4 5014 pch l=0.04u w=0.4u
m24156 5014 4389 4 5014 pch l=0.04u w=0.4u
m24157 VDDPOST 5747 5751 VDDPOST pch l=0.04u w=0.8u
m24158 VDDPOST 5869 5752 VDDPOST pch l=0.04u w=0.8u
m24159 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24160 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24161 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24162 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24163 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24164 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24165 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24166 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24167 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24168 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24169 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24170 5015 5014 5014 5014 pch l=0.04u w=0.4u
m24171 5765 4791 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24172 5708 5750 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24173 VDDPOST 4705 5765 VDDPOST pch l=0.04u w=0.8u
m24174 5766 5728 5751 VDDPOST pch l=0.04u w=0.8u
m24175 5767 5752 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24176 VDDPOST 5797 5708 VDDPOST pch l=0.04u w=0.8u
m24177 59591 5525 5766 VDDPOST pch l=0.04u w=0.24u
m24178 VDDPOST 5752 5767 VDDPOST pch l=0.04u w=0.8u
m24179 VDDPOST 5794 59591 VDDPOST pch l=0.04u w=0.24u
m24180 5768 5749 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24181 5770 5257 5750 VDDPOST pch l=0.04u w=0.8u
m24182 5772 5766 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24183 VDDPOST 5730 5768 VDDPOST pch l=0.04u w=0.8u
m24184 5773 5836 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24185 59853 5277 5770 VDDPOST pch l=0.04u w=0.12u
m24186 5783 5792 5771 VDDREF pch l=0.1u w=1u
m24187 VDDPOST 5790 59853 VDDPOST pch l=0.04u w=0.12u
m24188 5787 5627 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24189 5788 5768 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24190 5771 5792 5783 VDDREF pch l=0.1u w=1u
m24191 5789 POSTDIV1[0] VDDPOST VDDPOST pch l=0.04u w=0.12u
m24192 5790 5770 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24193 VDDPOST 5772 5787 VDDPOST pch l=0.04u w=0.8u
m24194 VDDPOST 5765 5788 VDDPOST pch l=0.04u w=0.8u
m24195 VDDPOST 5773 5789 VDDPOST pch l=0.04u w=0.4u
m24196 5788 5765 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24197 5789 5773 VDDPOST VDDPOST pch l=0.04u w=0.4u
m24198 5793 5277 5790 VDDPOST pch l=0.04u w=0.8u
m24199 VDDPOST 5768 5788 VDDPOST pch l=0.04u w=0.8u
m24200 5794 5787 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24201 60373 5792 5792 VDDREF pch l=0.25u w=1u
m24202 60497 5257 5793 VDDPOST pch l=0.04u w=0.12u
m24203 5795 5789 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24204 VDDPOST 5797 60497 VDDPOST pch l=0.04u w=0.12u
m24205 VDDREF 5792 60373 VDDREF pch l=0.25u w=1u
m24206 5796 BYPASS VDDPOST VDDPOST pch l=0.04u w=0.8u
m24207 VDDPOST 5824 5795 VDDPOST pch l=0.04u w=0.8u
m24208 5797 5793 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24209 VDDPOST 4953 5627 VDDPOST pch l=0.04u w=0.8u
m24210 60861 5783 VDDREF VDDREF pch l=0.25u w=1u
m24211 5799 5796 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24212 VDDPOST 5824 5798 VDDPOST pch l=0.04u w=0.8u
m24213 VDDPOST PD 5799 VDDPOST pch l=0.04u w=0.8u
m24214 5801 5790 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24215 5802 FOUT1PH0 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24216 5798 5807 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24217 5771 5783 60861 VDDREF pch l=0.25u w=1u
m24218 VDDPOST FOUT1PH0 5802 VDDPOST pch l=0.04u w=0.8u
m24219 VDDPOST 4933 5798 VDDPOST pch l=0.04u w=0.8u
m24220 5805 5799 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24221 5806 5797 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24222 5802 FOUT1PH0 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24223 61348 5783 5771 VDDREF pch l=0.25u w=1u
m24224 VDDPOST 4703 5805 VDDPOST pch l=0.04u w=0.8u
m24225 VDDPOST 5801 5806 VDDPOST pch l=0.04u w=0.8u
m24226 VDDPOST FOUT1PH0 5802 VDDPOST pch l=0.04u w=0.8u
m24227 VDDPOST 5831 5807 VDDPOST pch l=0.04u w=0.4u
m24228 VDDREF 5783 61348 VDDREF pch l=0.25u w=1u
m24229 5807 5831 VDDPOST VDDPOST pch l=0.04u w=0.4u
m24230 VDDPOST 5788 5811 VDDPOST pch l=0.04u w=0.8u
m24231 VDDPOST 5806 5812 VDDPOST pch l=0.04u w=0.8u
m24232 VDDPOST 5363 5813 VDDPOST pch l=0.04u w=0.8u
m24233 VDDPOST POSTDIV1[0] 5807 VDDPOST pch l=0.04u w=0.12u
m24234 61596 5783 VDDREF VDDREF pch l=0.25u w=1u
m24235 5817 5811 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24236 5818 5812 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24237 5819 5813 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24238 5771 5783 61596 VDDREF pch l=0.25u w=1u
m24239 5825 5901 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24240 5826 5902 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24241 5827 5903 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24242 VDDPOST 5829 5824 VDDPOST pch l=0.04u w=0.8u
m24243 VDDPOST 5788 5825 VDDPOST pch l=0.04u w=0.8u
m24244 VDDPOST 5806 5826 VDDPOST pch l=0.04u w=0.8u
m24245 VDDPOST 5363 5827 VDDPOST pch l=0.04u w=0.8u
m24246 61980 5824 VDDPOST VDDPOST pch l=0.04u w=0.12u
m24247 61981 5783 5771 VDDREF pch l=0.25u w=1u
m24248 5825 5788 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24249 5826 5806 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24250 5827 5363 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24251 5829 5864 61980 VDDPOST pch l=0.04u w=0.12u
m24252 VDDREF 5783 61981 VDDREF pch l=0.25u w=1u
m24253 5831 5837 5829 VDDPOST pch l=0.04u w=0.8u
m24254 FOUTPOSTDIV 5825 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24255 FOUT3 5826 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24256 FOUT1PH0 5827 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24257 VDDPOST 5825 FOUTPOSTDIV VDDPOST pch l=0.04u w=0.8u
m24258 VDDPOST 5826 FOUT3 VDDPOST pch l=0.04u w=0.8u
m24259 VDDPOST 5827 FOUT1PH0 VDDPOST pch l=0.04u w=0.8u
m24260 VDDPOST 5835 5831 VDDPOST pch l=0.04u w=0.8u
m24261 5783 5792 5771 VDDREF pch l=0.1u w=1u
m24262 FOUTPOSTDIV 5825 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24263 FOUT3 5826 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24264 FOUT1PH0 5827 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24265 62547 5831 VDDPOST VDDPOST pch l=0.04u w=0.12u
m24266 5771 5792 5783 VDDREF pch l=0.1u w=1u
m24267 VDDPOST 5825 FOUTPOSTDIV VDDPOST pch l=0.04u w=0.8u
m24268 VDDPOST 5826 FOUT3 VDDPOST pch l=0.04u w=0.8u
m24269 VDDPOST 5827 FOUT1PH0 VDDPOST pch l=0.04u w=0.8u
m24270 5835 5837 62547 VDDPOST pch l=0.04u w=0.12u
m24271 FOUTPOSTDIV 5825 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24272 FOUT3 5826 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24273 FOUT1PH0 5827 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24274 5836 5864 5835 VDDPOST pch l=0.04u w=0.8u
m24275 VDDPOST 5825 FOUTPOSTDIV VDDPOST pch l=0.04u w=0.8u
m24276 VDDPOST 5826 FOUT3 VDDPOST pch l=0.04u w=0.8u
m24277 VDDPOST 5827 FOUT1PH0 VDDPOST pch l=0.04u w=0.8u
m24278 FOUTPOSTDIV 5825 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24279 FOUT3 5826 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24280 FOUT1PH0 5827 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24281 VDDPOST 5864 5837 VDDPOST pch l=0.04u w=0.8u
m24282 VDDPOST 5825 FOUTPOSTDIV VDDPOST pch l=0.04u w=0.8u
m24283 VDDPOST 5826 FOUT3 VDDPOST pch l=0.04u w=0.8u
m24284 VDDPOST 5827 FOUT1PH0 VDDPOST pch l=0.04u w=0.8u
m24285 VDDPOST 5844 5836 VDDPOST pch l=0.04u w=0.8u
m24286 VDDPOST 5817 5838 VDDPOST pch l=0.04u w=0.8u
m24287 VDDPOST 5818 5839 VDDPOST pch l=0.04u w=0.8u
m24288 VDDPOST 5819 5840 VDDPOST pch l=0.04u w=0.8u
m24289 63464 5836 VDDPOST VDDPOST pch l=0.04u w=0.12u
m24290 5844 5864 63464 VDDPOST pch l=0.04u w=0.12u
m24291 5845 5817 5841 VDDPOST pch l=0.04u w=0.8u
m24292 5846 5818 5842 VDDPOST pch l=0.04u w=0.8u
m24293 5847 5819 5843 VDDPOST pch l=0.04u w=0.8u
m24294 5848 5859 5844 VDDPOST pch l=0.04u w=0.8u
m24295 63655 5838 5845 VDDPOST pch l=0.04u w=0.12u
m24296 63656 5839 5846 VDDPOST pch l=0.04u w=0.12u
m24297 63657 5840 5847 VDDPOST pch l=0.04u w=0.12u
m24298 VDDPOST 5849 63655 VDDPOST pch l=0.04u w=0.12u
m24299 VDDPOST 5850 63656 VDDPOST pch l=0.04u w=0.12u
m24300 VDDPOST 5851 63657 VDDPOST pch l=0.04u w=0.12u
m24301 VDDPOST 5853 5848 VDDPOST pch l=0.04u w=0.8u
m24302 5849 5841 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24303 5850 5842 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24304 5851 5843 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24305 63766 5848 VDDPOST VDDPOST pch l=0.04u w=0.12u
m24306 VDDPOST 5845 5849 VDDPOST pch l=0.04u w=0.8u
m24307 VDDPOST 5846 5850 VDDPOST pch l=0.04u w=0.8u
m24308 VDDPOST 5847 5851 VDDPOST pch l=0.04u w=0.8u
m24309 5853 5859 63766 VDDPOST pch l=0.04u w=0.12u
m24310 5795 5864 5853 VDDPOST pch l=0.04u w=0.8u
m24311 5855 5838 5849 VDDPOST pch l=0.04u w=0.8u
m24312 5856 5839 5850 VDDPOST pch l=0.04u w=0.8u
m24313 5857 5840 5851 VDDPOST pch l=0.04u w=0.8u
m24314 63900 5817 5855 VDDPOST pch l=0.04u w=0.24u
m24315 63901 5818 5856 VDDPOST pch l=0.04u w=0.24u
m24316 63902 5819 5857 VDDPOST pch l=0.04u w=0.24u
m24317 VDDPOST 5864 5859 VDDPOST pch l=0.04u w=0.8u
m24318 VDDPOST 5870 63900 VDDPOST pch l=0.04u w=0.24u
m24319 VDDPOST 5871 63901 VDDPOST pch l=0.04u w=0.24u
m24320 VDDPOST 5872 63902 VDDPOST pch l=0.04u w=0.24u
m24321 5861 5855 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24322 5862 5856 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24323 5863 5857 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24324 VDDPOST 4708 5864 VDDPOST pch l=0.04u w=0.8u
m24325 5866 5841 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24326 5867 5842 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24327 5868 5843 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24328 5864 4708 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24329 VDDPOST 5861 5866 VDDPOST pch l=0.04u w=0.8u
m24330 VDDPOST 5862 5867 VDDPOST pch l=0.04u w=0.8u
m24331 VDDPOST 5863 5868 VDDPOST pch l=0.04u w=0.8u
m24332 VDDPOST 4933 5864 VDDPOST pch l=0.04u w=0.8u
m24333 5870 5866 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24334 5871 5867 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24335 5872 5868 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24336 VDDPOST 5877 5869 VDDPOST pch l=0.04u w=0.4u
m24337 5869 5877 VDDPOST VDDPOST pch l=0.04u w=0.4u
m24338 VDDPOST 5817 5874 VDDPOST pch l=0.04u w=0.8u
m24339 VDDPOST 5818 5875 VDDPOST pch l=0.04u w=0.8u
m24340 VDDPOST 5819 5876 VDDPOST pch l=0.04u w=0.8u
m24341 VDDPOST 4925 5869 VDDPOST pch l=0.04u w=0.12u
m24342 5878 5817 5870 VDDPOST pch l=0.04u w=0.8u
m24343 5879 5818 5871 VDDPOST pch l=0.04u w=0.8u
m24344 5880 5819 5872 VDDPOST pch l=0.04u w=0.8u
m24345 VDDPOST 5881 5877 VDDPOST pch l=0.04u w=0.8u
m24346 64738 5874 5878 VDDPOST pch l=0.04u w=0.12u
m24347 64739 5875 5879 VDDPOST pch l=0.04u w=0.12u
m24348 64740 5876 5880 VDDPOST pch l=0.04u w=0.12u
m24349 64742 5877 VDDPOST VDDPOST pch l=0.04u w=0.12u
m24350 VDDPOST 5883 64738 VDDPOST pch l=0.04u w=0.12u
m24351 VDDPOST 5884 64739 VDDPOST pch l=0.04u w=0.12u
m24352 VDDPOST 5885 64740 VDDPOST pch l=0.04u w=0.12u
m24353 5881 5899 64742 VDDPOST pch l=0.04u w=0.12u
m24354 5883 5841 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24355 5884 5842 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24356 5885 5843 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24357 5886 5895 5881 VDDPOST pch l=0.04u w=0.8u
m24358 VDDPOST 5878 5883 VDDPOST pch l=0.04u w=0.8u
m24359 VDDPOST 5879 5884 VDDPOST pch l=0.04u w=0.8u
m24360 VDDPOST 5880 5885 VDDPOST pch l=0.04u w=0.8u
m24361 VDDPOST 5890 5886 VDDPOST pch l=0.04u w=0.8u
m24362 5887 5874 5883 VDDPOST pch l=0.04u w=0.8u
m24363 5888 5875 5884 VDDPOST pch l=0.04u w=0.8u
m24364 5889 5876 5885 VDDPOST pch l=0.04u w=0.8u
m24365 65103 5886 VDDPOST VDDPOST pch l=0.04u w=0.12u
m24366 65326 5817 5887 VDDPOST pch l=0.04u w=0.24u
m24367 65327 5818 5888 VDDPOST pch l=0.04u w=0.24u
m24368 65328 5819 5889 VDDPOST pch l=0.04u w=0.24u
m24369 5890 5895 65103 VDDPOST pch l=0.04u w=0.12u
m24370 VDDPOST 5901 65326 VDDPOST pch l=0.04u w=0.24u
m24371 VDDPOST 5902 65327 VDDPOST pch l=0.04u w=0.24u
m24372 VDDPOST 5903 65328 VDDPOST pch l=0.04u w=0.24u
m24373 5891 5899 5890 VDDPOST pch l=0.04u w=0.8u
m24374 5892 5887 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24375 5893 5888 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24376 5894 5889 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24377 VDDPOST 5899 5895 VDDPOST pch l=0.04u w=0.8u
m24378 5896 5841 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24379 5897 5842 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24380 5898 5843 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24381 VDDPOST 5892 5896 VDDPOST pch l=0.04u w=0.8u
m24382 VDDPOST 5893 5897 VDDPOST pch l=0.04u w=0.8u
m24383 VDDPOST 5894 5898 VDDPOST pch l=0.04u w=0.8u
m24384 VDDPOST 4708 5899 VDDPOST pch l=0.04u w=0.4u
m24385 5901 5896 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24386 5902 5897 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24387 5903 5898 VDDPOST VDDPOST pch l=0.04u w=0.8u
m24388 5899 4708 VDDPOST VDDPOST pch l=0.04u w=0.4u
m24389 VDDPOST 4925 5899 VDDPOST pch l=0.04u w=0.12u
m24390 VDDPOST 5877 5891 VDDPOST pch l=0.04u w=0.8u
m24391 VDDPOST 5805 5841 VDDPOST pch l=0.04u w=0.8u
m24392 VDDPOST 4953 5842 VDDPOST pch l=0.04u w=0.8u
m24393 VDDPOST 4953 5843 VDDPOST pch l=0.04u w=0.8u
x24394 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24395 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24396 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24397 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24398 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24399 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24400 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24401 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24402 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24403 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24404 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24405 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24406 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24407 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24408 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24409 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24410 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24411 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24412 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24413 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24414 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24415 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24416 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24417 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24418 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24419 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24420 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24421 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24422 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24423 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24424 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24425 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24426 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24427 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24428 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24429 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24430 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24431 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24432 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24433 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24434 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24435 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24436 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24437 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24438 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24439 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24440 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24441 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24442 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24443 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24444 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24445 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24446 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24447 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24448 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24449 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24450 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24451 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24452 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24453 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24454 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24455 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24456 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24457 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24458 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24459 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24460 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24461 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24462 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24463 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24464 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24465 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24466 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24467 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24468 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24469 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24470 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24471 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24472 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24473 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24474 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24475 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24476 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24477 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24478 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24479 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24480 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24481 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24482 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24483 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24484 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24485 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24486 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24487 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24488 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24489 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24490 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24491 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24492 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24493 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24494 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24495 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24496 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24497 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24498 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24499 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24500 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24501 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24502 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24503 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24504 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24505 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24506 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24507 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24508 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24509 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24510 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24511 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24512 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24513 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24514 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24515 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24516 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24517 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24518 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24519 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24520 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24521 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24522 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24523 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24524 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24525 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24526 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24527 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24528 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24529 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24530 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24531 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24532 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24533 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24534 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24535 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24536 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24537 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24538 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24539 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24540 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24541 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24542 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24543 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24544 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24545 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24546 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24547 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24548 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24549 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24550 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24551 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24552 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24553 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24554 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24555 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24556 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24557 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24558 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24559 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24560 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24561 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24562 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24563 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24564 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24565 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24566 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24567 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24568 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24569 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24570 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24571 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24572 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24573 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24574 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24575 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24576 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24577 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24578 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24579 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24580 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24581 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24582 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24583 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24584 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24585 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24586 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24587 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24588 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24589 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24590 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24591 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24592 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24593 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24594 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24595 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24596 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24597 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24598 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24599 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24600 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24601 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24602 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24603 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24604 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24605 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24606 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24607 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24608 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24609 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24610 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24611 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24612 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24613 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24614 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24615 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24616 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24617 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24618 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24619 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24620 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24621 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24622 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24623 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24624 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24625 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24626 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24627 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24628 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24629 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24630 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24631 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24632 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24633 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24634 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24635 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24636 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24637 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24638 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24639 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24640 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24641 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24642 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24643 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24644 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24645 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24646 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24647 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24648 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24649 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24650 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24651 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24652 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24653 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24654 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24655 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24656 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24657 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24658 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24659 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24660 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24661 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24662 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24663 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24664 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24665 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24666 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24667 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24668 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24669 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24670 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24671 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24672 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24673 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24674 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24675 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24676 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24677 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24678 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24679 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24680 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24681 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24682 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24683 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24684 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24685 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24686 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24687 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24688 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24689 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24690 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24691 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24692 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24693 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24694 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24695 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24696 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24697 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24698 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24699 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24700 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24701 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24702 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24703 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24704 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24705 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24706 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24707 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24708 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24709 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24710 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24711 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24712 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24713 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24714 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24715 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24716 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24717 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24718 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24719 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24720 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24721 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24722 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24723 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24724 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24725 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24726 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24727 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24728 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24729 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24730 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24731 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24732 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24733 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24734 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24735 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24736 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24737 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24738 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24739 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24740 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24741 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24742 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24743 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24744 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24745 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24746 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24747 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24748 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24749 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24750 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24751 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24752 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24753 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24754 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24755 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24756 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24757 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24758 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24759 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24760 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24761 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24762 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24763 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24764 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24765 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24766 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24767 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24768 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24769 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24770 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24771 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24772 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24773 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24774 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24775 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24776 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24777 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24778 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24779 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24780 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24781 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24782 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24783 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24784 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24785 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24786 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24787 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24788 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24789 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24790 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24791 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24792 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24793 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24794 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24795 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24796 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24797 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24798 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24799 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24800 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24801 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24802 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24803 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24804 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24805 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24806 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24807 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24808 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24809 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24810 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24811 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24812 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24813 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24814 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24815 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24816 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24817 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24818 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24819 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24820 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24821 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24822 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24823 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24824 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24825 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24826 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24827 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24828 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24829 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24830 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24831 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24832 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24833 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24834 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24835 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24836 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24837 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24838 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24839 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24840 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24841 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24842 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24843 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24844 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24845 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24846 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24847 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24848 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24849 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24850 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24851 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24852 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24853 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24854 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24855 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24856 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24857 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24858 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24859 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24860 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24861 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24862 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24863 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24864 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24865 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24866 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24867 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24868 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24869 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24870 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24871 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24872 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24873 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24874 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24875 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24876 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24877 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24878 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24879 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24880 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24881 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24882 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24883 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24884 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24885 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24886 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24887 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24888 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24889 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24890 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24891 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24892 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24893 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24894 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24895 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24896 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24897 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24898 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24899 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24900 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24901 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24902 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24903 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24904 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24905 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24906 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24907 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24908 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24909 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24910 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24911 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24912 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24913 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24914 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24915 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24916 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24917 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24918 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24919 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24920 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24921 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24922 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24923 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24924 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24925 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24926 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24927 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24928 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24929 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24930 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24931 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24932 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24933 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24934 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24935 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24936 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24937 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24938 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24939 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24940 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24941 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24942 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24943 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24944 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24945 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24946 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24947 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24948 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24949 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24950 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24951 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24952 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24953 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24954 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24955 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24956 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24957 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24958 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24959 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24960 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24961 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24962 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24963 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24964 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24965 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24966 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24967 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24968 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24969 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24970 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24971 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24972 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24973 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24974 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24975 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24976 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24977 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24978 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24979 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24980 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24981 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24982 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24983 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24984 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24985 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24986 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24987 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24988 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x24989 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24990 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24991 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24992 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24993 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24994 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24995 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24996 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24997 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24998 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x24999 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25000 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25001 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25002 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25003 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25004 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25005 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25006 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25007 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25008 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25009 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25010 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25011 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25012 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25013 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25014 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25015 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25016 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25017 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25018 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25019 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25020 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25021 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25022 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25023 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25024 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25025 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25026 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25027 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25028 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25029 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25030 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25031 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25032 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25033 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25034 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25035 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25036 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25037 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25038 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25039 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25040 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25041 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25042 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25043 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25044 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25045 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25046 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25047 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25048 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25049 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25050 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25051 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25052 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25053 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25054 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25055 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25056 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25057 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25058 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25059 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25060 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25061 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25062 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25063 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25064 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25065 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25066 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25067 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25068 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25069 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25070 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25071 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25072 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25073 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25074 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25075 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25076 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25077 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25078 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25079 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25080 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25081 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25082 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25083 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25084 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25085 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25086 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25087 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25088 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25089 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25090 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25091 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25092 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25093 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25094 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25095 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25096 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25097 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25098 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25099 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25100 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25101 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25102 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25103 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25104 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25105 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25106 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25107 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25108 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25109 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25110 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25111 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25112 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25113 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25114 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25115 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25116 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25117 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25118 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25119 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25120 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25121 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25122 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25123 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25124 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25125 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25126 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25127 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25128 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25129 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25130 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25131 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25132 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25133 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25134 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25135 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25136 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25137 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25138 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25139 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25140 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25141 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25142 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25143 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25144 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25145 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25146 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25147 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25148 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25149 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25150 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25151 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25152 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25153 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25154 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25155 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25156 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25157 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25158 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25159 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25160 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25161 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25162 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25163 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25164 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25165 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25166 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25167 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25168 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25169 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25170 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25171 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25172 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25173 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25174 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25175 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25176 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25177 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25178 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25179 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25180 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25181 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25182 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25183 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25184 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25185 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25186 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25187 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25188 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25189 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25190 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25191 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25192 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25193 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25194 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25195 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25196 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25197 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25198 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25199 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25200 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25201 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25202 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25203 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25204 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25205 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25206 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25207 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25208 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25209 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25210 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25211 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25212 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25213 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25214 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25215 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25216 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25217 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25218 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25219 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25220 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25221 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25222 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25223 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25224 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25225 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25226 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25227 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25228 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25229 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25230 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25231 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25232 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25233 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25234 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25235 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25236 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25237 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25238 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25239 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25240 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25241 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25242 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25243 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25244 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25245 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25246 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25247 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25248 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25249 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25250 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25251 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25252 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25253 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25254 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25255 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25256 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25257 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25258 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25259 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25260 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25261 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25262 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25263 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25264 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25265 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25266 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25267 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25268 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25269 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25270 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25271 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25272 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25273 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25274 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25275 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25276 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25277 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25278 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25279 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25280 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25281 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25282 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25283 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25284 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25285 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25286 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25287 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25288 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25289 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25290 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25291 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25292 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25293 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25294 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25295 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25296 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25297 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25298 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25299 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25300 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25301 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25302 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25303 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25304 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25305 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25306 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25307 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25308 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25309 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25310 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25311 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25312 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25313 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25314 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25315 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25316 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25317 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25318 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25319 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25320 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25321 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25322 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25323 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25324 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25325 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25326 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25327 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25328 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25329 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25330 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25331 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25332 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25333 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25334 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25335 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25336 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25337 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25338 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25339 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25340 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25341 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25342 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25343 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25344 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25345 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25346 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25347 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25348 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25349 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25350 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25351 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25352 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25353 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25354 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25355 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25356 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25357 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25358 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25359 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25360 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25361 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25362 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25363 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25364 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25365 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25366 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25367 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25368 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25369 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25370 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25371 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25372 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25373 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25374 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25375 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25376 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25377 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25378 VDDPOST VSS nmoscap_18 lr=1.9u wr=2.98u
x25379 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25380 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25381 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25382 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25383 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25384 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25385 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25386 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25387 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25388 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25389 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25390 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25391 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25392 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25393 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25394 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25395 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25396 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25397 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25398 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25399 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25400 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25401 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25402 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25403 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25404 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25405 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25406 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25407 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25408 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25409 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25410 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25411 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25412 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25413 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25414 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25415 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25416 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25417 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25418 4 VSS nmoscap_18 lr=1.9u wr=2.98u
x25419 5528 5339 nmoscap_18 lr=2.1u wr=2.4u
x25420 5528 5339 nmoscap_18 lr=2.1u wr=2.4u
x25421 5528 5339 nmoscap_18 lr=2.1u wr=2.4u
x25422 5528 5339 nmoscap_18 lr=2.1u wr=2.4u
x25423 5528 5339 nmoscap_18 lr=2.1u wr=2.4u
x25424 5528 5339 nmoscap_18 lr=2.1u wr=2.4u
x25425 5339 5528 nmoscap_18 lr=2.1u wr=2.4u
x25426 5339 5528 nmoscap_18 lr=2.1u wr=2.4u
x25427 5339 5528 nmoscap_18 lr=2.1u wr=2.4u
x25428 5339 5528 nmoscap_18 lr=2.1u wr=2.4u
x25429 5339 5528 nmoscap_18 lr=2.1u wr=2.4u
x25430 5339 5528 nmoscap_18 lr=2.1u wr=2.4u
.ends PLLTS40GFRAC
